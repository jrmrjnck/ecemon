module Protag_Fight
(
   input            clock, 
   input      [7:0] x,
   input      [7:0] y, 
   input      [7:0] loc_x, 
   input      [7:0] loc_y, 
   output reg       on,
   output reg [1:0] color
);

   localparam WIDTH = 8'd64,
              HEIGHT = 8'd64;

   // Buffer the scan coordinates to synchronize
   // with the ROM data output
   always @( posedge clock ) begin
    on <= (x >= loc_x && x <= (loc_x+(WIDTH-1)))
          && (y >= loc_y && y <= (loc_y+(HEIGHT-1)));
   end

   reg [11:0] addr;
   always @( posedge clock )
      addr <= {y[5:0]-loc_y[5:0],x[5:0]-loc_x[5:0]};

always @(*) begin
   case( addr )
      12'h000: color = 2'b11;
      12'h001: color = 2'b11;
      12'h002: color = 2'b11;
      12'h003: color = 2'b11;
      12'h004: color = 2'b11;
      12'h005: color = 2'b11;
      12'h006: color = 2'b11;
      12'h007: color = 2'b11;
      12'h008: color = 2'b11;
      12'h009: color = 2'b11;
      12'h00a: color = 2'b11;
      12'h00b: color = 2'b11;
      12'h00c: color = 2'b11;
      12'h00d: color = 2'b11;
      12'h00e: color = 2'b11;
      12'h00f: color = 2'b11;
      12'h010: color = 2'b11;
      12'h011: color = 2'b11;
      12'h012: color = 2'b11;
      12'h013: color = 2'b11;
      12'h014: color = 2'b11;
      12'h015: color = 2'b11;
      12'h016: color = 2'b11;
      12'h017: color = 2'b11;
      12'h018: color = 2'b11;
      12'h019: color = 2'b11;
      12'h01a: color = 2'b11;
      12'h01b: color = 2'b11;
      12'h01c: color = 2'b11;
      12'h01d: color = 2'b11;
      12'h01e: color = 2'b00;
      12'h01f: color = 2'b00;
      12'h020: color = 2'b00;
      12'h021: color = 2'b00;
      12'h022: color = 2'b00;
      12'h023: color = 2'b00;
      12'h024: color = 2'b00;
      12'h025: color = 2'b01;
      12'h026: color = 2'b01;
      12'h027: color = 2'b11;
      12'h028: color = 2'b11;
      12'h029: color = 2'b11;
      12'h02a: color = 2'b11;
      12'h02b: color = 2'b11;
      12'h02c: color = 2'b11;
      12'h02d: color = 2'b11;
      12'h02e: color = 2'b11;
      12'h02f: color = 2'b11;
      12'h030: color = 2'b11;
      12'h031: color = 2'b11;
      12'h032: color = 2'b11;
      12'h033: color = 2'b11;
      12'h034: color = 2'b11;
      12'h035: color = 2'b11;
      12'h036: color = 2'b11;
      12'h037: color = 2'b11;
      12'h038: color = 2'b11;
      12'h039: color = 2'b11;
      12'h03a: color = 2'b11;
      12'h03b: color = 2'b11;
      12'h03c: color = 2'b11;
      12'h03d: color = 2'b11;
      12'h03e: color = 2'b11;
      12'h03f: color = 2'b11;
      12'h040: color = 2'b11;
      12'h041: color = 2'b11;
      12'h042: color = 2'b11;
      12'h043: color = 2'b11;
      12'h044: color = 2'b11;
      12'h045: color = 2'b11;
      12'h046: color = 2'b11;
      12'h047: color = 2'b11;
      12'h048: color = 2'b11;
      12'h049: color = 2'b11;
      12'h04a: color = 2'b11;
      12'h04b: color = 2'b11;
      12'h04c: color = 2'b11;
      12'h04d: color = 2'b11;
      12'h04e: color = 2'b11;
      12'h04f: color = 2'b11;
      12'h050: color = 2'b11;
      12'h051: color = 2'b11;
      12'h052: color = 2'b11;
      12'h053: color = 2'b11;
      12'h054: color = 2'b11;
      12'h055: color = 2'b11;
      12'h056: color = 2'b11;
      12'h057: color = 2'b11;
      12'h058: color = 2'b11;
      12'h059: color = 2'b11;
      12'h05a: color = 2'b11;
      12'h05b: color = 2'b11;
      12'h05c: color = 2'b11;
      12'h05d: color = 2'b11;
      12'h05e: color = 2'b00;
      12'h05f: color = 2'b00;
      12'h060: color = 2'b00;
      12'h061: color = 2'b00;
      12'h062: color = 2'b00;
      12'h063: color = 2'b00;
      12'h064: color = 2'b00;
      12'h065: color = 2'b01;
      12'h066: color = 2'b01;
      12'h067: color = 2'b11;
      12'h068: color = 2'b11;
      12'h069: color = 2'b11;
      12'h06a: color = 2'b11;
      12'h06b: color = 2'b11;
      12'h06c: color = 2'b11;
      12'h06d: color = 2'b11;
      12'h06e: color = 2'b11;
      12'h06f: color = 2'b11;
      12'h070: color = 2'b11;
      12'h071: color = 2'b11;
      12'h072: color = 2'b11;
      12'h073: color = 2'b11;
      12'h074: color = 2'b11;
      12'h075: color = 2'b11;
      12'h076: color = 2'b11;
      12'h077: color = 2'b11;
      12'h078: color = 2'b11;
      12'h079: color = 2'b11;
      12'h07a: color = 2'b11;
      12'h07b: color = 2'b11;
      12'h07c: color = 2'b11;
      12'h07d: color = 2'b11;
      12'h07e: color = 2'b11;
      12'h07f: color = 2'b11;
      12'h080: color = 2'b11;
      12'h081: color = 2'b11;
      12'h082: color = 2'b11;
      12'h083: color = 2'b11;
      12'h084: color = 2'b11;
      12'h085: color = 2'b11;
      12'h086: color = 2'b11;
      12'h087: color = 2'b11;
      12'h088: color = 2'b11;
      12'h089: color = 2'b11;
      12'h08a: color = 2'b11;
      12'h08b: color = 2'b11;
      12'h08c: color = 2'b11;
      12'h08d: color = 2'b11;
      12'h08e: color = 2'b11;
      12'h08f: color = 2'b11;
      12'h090: color = 2'b11;
      12'h091: color = 2'b11;
      12'h092: color = 2'b11;
      12'h093: color = 2'b11;
      12'h094: color = 2'b11;
      12'h095: color = 2'b11;
      12'h096: color = 2'b11;
      12'h097: color = 2'b11;
      12'h098: color = 2'b11;
      12'h099: color = 2'b00;
      12'h09a: color = 2'b00;
      12'h09b: color = 2'b00;
      12'h09c: color = 2'b00;
      12'h09d: color = 2'b00;
      12'h09e: color = 2'b10;
      12'h09f: color = 2'b10;
      12'h0a0: color = 2'b10;
      12'h0a1: color = 2'b10;
      12'h0a2: color = 2'b10;
      12'h0a3: color = 2'b10;
      12'h0a4: color = 2'b10;
      12'h0a5: color = 2'b10;
      12'h0a6: color = 2'b10;
      12'h0a7: color = 2'b00;
      12'h0a8: color = 2'b00;
      12'h0a9: color = 2'b00;
      12'h0aa: color = 2'b00;
      12'h0ab: color = 2'b11;
      12'h0ac: color = 2'b11;
      12'h0ad: color = 2'b11;
      12'h0ae: color = 2'b11;
      12'h0af: color = 2'b11;
      12'h0b0: color = 2'b11;
      12'h0b1: color = 2'b11;
      12'h0b2: color = 2'b11;
      12'h0b3: color = 2'b11;
      12'h0b4: color = 2'b11;
      12'h0b5: color = 2'b11;
      12'h0b6: color = 2'b11;
      12'h0b7: color = 2'b11;
      12'h0b8: color = 2'b11;
      12'h0b9: color = 2'b11;
      12'h0ba: color = 2'b11;
      12'h0bb: color = 2'b11;
      12'h0bc: color = 2'b11;
      12'h0bd: color = 2'b11;
      12'h0be: color = 2'b11;
      12'h0bf: color = 2'b11;
      12'h0c0: color = 2'b11;
      12'h0c1: color = 2'b11;
      12'h0c2: color = 2'b11;
      12'h0c3: color = 2'b11;
      12'h0c4: color = 2'b11;
      12'h0c5: color = 2'b11;
      12'h0c6: color = 2'b11;
      12'h0c7: color = 2'b11;
      12'h0c8: color = 2'b11;
      12'h0c9: color = 2'b11;
      12'h0ca: color = 2'b11;
      12'h0cb: color = 2'b11;
      12'h0cc: color = 2'b11;
      12'h0cd: color = 2'b11;
      12'h0ce: color = 2'b11;
      12'h0cf: color = 2'b11;
      12'h0d0: color = 2'b11;
      12'h0d1: color = 2'b11;
      12'h0d2: color = 2'b11;
      12'h0d3: color = 2'b11;
      12'h0d4: color = 2'b11;
      12'h0d5: color = 2'b11;
      12'h0d6: color = 2'b11;
      12'h0d7: color = 2'b11;
      12'h0d8: color = 2'b11;
      12'h0d9: color = 2'b00;
      12'h0da: color = 2'b00;
      12'h0db: color = 2'b00;
      12'h0dc: color = 2'b00;
      12'h0dd: color = 2'b00;
      12'h0de: color = 2'b10;
      12'h0df: color = 2'b10;
      12'h0e0: color = 2'b10;
      12'h0e1: color = 2'b10;
      12'h0e2: color = 2'b10;
      12'h0e3: color = 2'b10;
      12'h0e4: color = 2'b10;
      12'h0e5: color = 2'b10;
      12'h0e6: color = 2'b10;
      12'h0e7: color = 2'b00;
      12'h0e8: color = 2'b00;
      12'h0e9: color = 2'b00;
      12'h0ea: color = 2'b00;
      12'h0eb: color = 2'b11;
      12'h0ec: color = 2'b11;
      12'h0ed: color = 2'b11;
      12'h0ee: color = 2'b11;
      12'h0ef: color = 2'b11;
      12'h0f0: color = 2'b11;
      12'h0f1: color = 2'b11;
      12'h0f2: color = 2'b11;
      12'h0f3: color = 2'b11;
      12'h0f4: color = 2'b11;
      12'h0f5: color = 2'b11;
      12'h0f6: color = 2'b11;
      12'h0f7: color = 2'b11;
      12'h0f8: color = 2'b11;
      12'h0f9: color = 2'b11;
      12'h0fa: color = 2'b11;
      12'h0fb: color = 2'b11;
      12'h0fc: color = 2'b11;
      12'h0fd: color = 2'b11;
      12'h0fe: color = 2'b11;
      12'h0ff: color = 2'b11;
      12'h100: color = 2'b11;
      12'h101: color = 2'b11;
      12'h102: color = 2'b11;
      12'h103: color = 2'b11;
      12'h104: color = 2'b11;
      12'h105: color = 2'b11;
      12'h106: color = 2'b11;
      12'h107: color = 2'b11;
      12'h108: color = 2'b11;
      12'h109: color = 2'b11;
      12'h10a: color = 2'b11;
      12'h10b: color = 2'b11;
      12'h10c: color = 2'b11;
      12'h10d: color = 2'b11;
      12'h10e: color = 2'b11;
      12'h10f: color = 2'b11;
      12'h110: color = 2'b11;
      12'h111: color = 2'b11;
      12'h112: color = 2'b11;
      12'h113: color = 2'b11;
      12'h114: color = 2'b11;
      12'h115: color = 2'b00;
      12'h116: color = 2'b00;
      12'h117: color = 2'b00;
      12'h118: color = 2'b00;
      12'h119: color = 2'b10;
      12'h11a: color = 2'b10;
      12'h11b: color = 2'b10;
      12'h11c: color = 2'b10;
      12'h11d: color = 2'b10;
      12'h11e: color = 2'b10;
      12'h11f: color = 2'b10;
      12'h120: color = 2'b10;
      12'h121: color = 2'b10;
      12'h122: color = 2'b10;
      12'h123: color = 2'b10;
      12'h124: color = 2'b10;
      12'h125: color = 2'b10;
      12'h126: color = 2'b10;
      12'h127: color = 2'b10;
      12'h128: color = 2'b10;
      12'h129: color = 2'b10;
      12'h12a: color = 2'b10;
      12'h12b: color = 2'b00;
      12'h12c: color = 2'b00;
      12'h12d: color = 2'b00;
      12'h12e: color = 2'b11;
      12'h12f: color = 2'b11;
      12'h130: color = 2'b11;
      12'h131: color = 2'b11;
      12'h132: color = 2'b11;
      12'h133: color = 2'b11;
      12'h134: color = 2'b11;
      12'h135: color = 2'b11;
      12'h136: color = 2'b11;
      12'h137: color = 2'b11;
      12'h138: color = 2'b11;
      12'h139: color = 2'b11;
      12'h13a: color = 2'b11;
      12'h13b: color = 2'b11;
      12'h13c: color = 2'b11;
      12'h13d: color = 2'b11;
      12'h13e: color = 2'b11;
      12'h13f: color = 2'b11;
      12'h140: color = 2'b11;
      12'h141: color = 2'b11;
      12'h142: color = 2'b11;
      12'h143: color = 2'b11;
      12'h144: color = 2'b11;
      12'h145: color = 2'b11;
      12'h146: color = 2'b11;
      12'h147: color = 2'b11;
      12'h148: color = 2'b11;
      12'h149: color = 2'b11;
      12'h14a: color = 2'b11;
      12'h14b: color = 2'b11;
      12'h14c: color = 2'b11;
      12'h14d: color = 2'b11;
      12'h14e: color = 2'b11;
      12'h14f: color = 2'b11;
      12'h150: color = 2'b11;
      12'h151: color = 2'b11;
      12'h152: color = 2'b11;
      12'h153: color = 2'b11;
      12'h154: color = 2'b11;
      12'h155: color = 2'b00;
      12'h156: color = 2'b00;
      12'h157: color = 2'b00;
      12'h158: color = 2'b00;
      12'h159: color = 2'b10;
      12'h15a: color = 2'b10;
      12'h15b: color = 2'b10;
      12'h15c: color = 2'b10;
      12'h15d: color = 2'b10;
      12'h15e: color = 2'b10;
      12'h15f: color = 2'b10;
      12'h160: color = 2'b10;
      12'h161: color = 2'b10;
      12'h162: color = 2'b10;
      12'h163: color = 2'b10;
      12'h164: color = 2'b10;
      12'h165: color = 2'b10;
      12'h166: color = 2'b10;
      12'h167: color = 2'b10;
      12'h168: color = 2'b10;
      12'h169: color = 2'b10;
      12'h16a: color = 2'b10;
      12'h16b: color = 2'b00;
      12'h16c: color = 2'b00;
      12'h16d: color = 2'b00;
      12'h16e: color = 2'b11;
      12'h16f: color = 2'b11;
      12'h170: color = 2'b11;
      12'h171: color = 2'b11;
      12'h172: color = 2'b11;
      12'h173: color = 2'b11;
      12'h174: color = 2'b11;
      12'h175: color = 2'b11;
      12'h176: color = 2'b11;
      12'h177: color = 2'b11;
      12'h178: color = 2'b11;
      12'h179: color = 2'b11;
      12'h17a: color = 2'b11;
      12'h17b: color = 2'b11;
      12'h17c: color = 2'b11;
      12'h17d: color = 2'b11;
      12'h17e: color = 2'b11;
      12'h17f: color = 2'b11;
      12'h180: color = 2'b11;
      12'h181: color = 2'b11;
      12'h182: color = 2'b11;
      12'h183: color = 2'b11;
      12'h184: color = 2'b11;
      12'h185: color = 2'b11;
      12'h186: color = 2'b11;
      12'h187: color = 2'b11;
      12'h188: color = 2'b11;
      12'h189: color = 2'b11;
      12'h18a: color = 2'b11;
      12'h18b: color = 2'b11;
      12'h18c: color = 2'b11;
      12'h18d: color = 2'b11;
      12'h18e: color = 2'b11;
      12'h18f: color = 2'b11;
      12'h190: color = 2'b00;
      12'h191: color = 2'b00;
      12'h192: color = 2'b00;
      12'h193: color = 2'b00;
      12'h194: color = 2'b00;
      12'h195: color = 2'b01;
      12'h196: color = 2'b01;
      12'h197: color = 2'b01;
      12'h198: color = 2'b01;
      12'h199: color = 2'b01;
      12'h19a: color = 2'b01;
      12'h19b: color = 2'b10;
      12'h19c: color = 2'b10;
      12'h19d: color = 2'b10;
      12'h19e: color = 2'b01;
      12'h19f: color = 2'b01;
      12'h1a0: color = 2'b10;
      12'h1a1: color = 2'b10;
      12'h1a2: color = 2'b10;
      12'h1a3: color = 2'b10;
      12'h1a4: color = 2'b10;
      12'h1a5: color = 2'b10;
      12'h1a6: color = 2'b10;
      12'h1a7: color = 2'b10;
      12'h1a8: color = 2'b10;
      12'h1a9: color = 2'b10;
      12'h1aa: color = 2'b10;
      12'h1ab: color = 2'b00;
      12'h1ac: color = 2'b00;
      12'h1ad: color = 2'b00;
      12'h1ae: color = 2'b11;
      12'h1af: color = 2'b11;
      12'h1b0: color = 2'b11;
      12'h1b1: color = 2'b11;
      12'h1b2: color = 2'b11;
      12'h1b3: color = 2'b11;
      12'h1b4: color = 2'b11;
      12'h1b5: color = 2'b11;
      12'h1b6: color = 2'b11;
      12'h1b7: color = 2'b11;
      12'h1b8: color = 2'b11;
      12'h1b9: color = 2'b11;
      12'h1ba: color = 2'b11;
      12'h1bb: color = 2'b11;
      12'h1bc: color = 2'b11;
      12'h1bd: color = 2'b11;
      12'h1be: color = 2'b11;
      12'h1bf: color = 2'b11;
      12'h1c0: color = 2'b11;
      12'h1c1: color = 2'b11;
      12'h1c2: color = 2'b11;
      12'h1c3: color = 2'b11;
      12'h1c4: color = 2'b11;
      12'h1c5: color = 2'b11;
      12'h1c6: color = 2'b11;
      12'h1c7: color = 2'b11;
      12'h1c8: color = 2'b11;
      12'h1c9: color = 2'b11;
      12'h1ca: color = 2'b11;
      12'h1cb: color = 2'b11;
      12'h1cc: color = 2'b11;
      12'h1cd: color = 2'b11;
      12'h1ce: color = 2'b11;
      12'h1cf: color = 2'b11;
      12'h1d0: color = 2'b00;
      12'h1d1: color = 2'b00;
      12'h1d2: color = 2'b00;
      12'h1d3: color = 2'b00;
      12'h1d4: color = 2'b00;
      12'h1d5: color = 2'b01;
      12'h1d6: color = 2'b01;
      12'h1d7: color = 2'b01;
      12'h1d8: color = 2'b01;
      12'h1d9: color = 2'b01;
      12'h1da: color = 2'b01;
      12'h1db: color = 2'b10;
      12'h1dc: color = 2'b10;
      12'h1dd: color = 2'b10;
      12'h1de: color = 2'b01;
      12'h1df: color = 2'b01;
      12'h1e0: color = 2'b10;
      12'h1e1: color = 2'b10;
      12'h1e2: color = 2'b10;
      12'h1e3: color = 2'b10;
      12'h1e4: color = 2'b10;
      12'h1e5: color = 2'b10;
      12'h1e6: color = 2'b10;
      12'h1e7: color = 2'b10;
      12'h1e8: color = 2'b10;
      12'h1e9: color = 2'b10;
      12'h1ea: color = 2'b10;
      12'h1eb: color = 2'b00;
      12'h1ec: color = 2'b00;
      12'h1ed: color = 2'b00;
      12'h1ee: color = 2'b11;
      12'h1ef: color = 2'b11;
      12'h1f0: color = 2'b11;
      12'h1f1: color = 2'b11;
      12'h1f2: color = 2'b11;
      12'h1f3: color = 2'b11;
      12'h1f4: color = 2'b11;
      12'h1f5: color = 2'b11;
      12'h1f6: color = 2'b11;
      12'h1f7: color = 2'b11;
      12'h1f8: color = 2'b11;
      12'h1f9: color = 2'b11;
      12'h1fa: color = 2'b11;
      12'h1fb: color = 2'b11;
      12'h1fc: color = 2'b11;
      12'h1fd: color = 2'b11;
      12'h1fe: color = 2'b11;
      12'h1ff: color = 2'b11;
      12'h200: color = 2'b11;
      12'h201: color = 2'b11;
      12'h202: color = 2'b11;
      12'h203: color = 2'b11;
      12'h204: color = 2'b11;
      12'h205: color = 2'b11;
      12'h206: color = 2'b11;
      12'h207: color = 2'b11;
      12'h208: color = 2'b11;
      12'h209: color = 2'b11;
      12'h20a: color = 2'b11;
      12'h20b: color = 2'b11;
      12'h20c: color = 2'b11;
      12'h20d: color = 2'b11;
      12'h20e: color = 2'b11;
      12'h20f: color = 2'b11;
      12'h210: color = 2'b00;
      12'h211: color = 2'b00;
      12'h212: color = 2'b00;
      12'h213: color = 2'b00;
      12'h214: color = 2'b00;
      12'h215: color = 2'b01;
      12'h216: color = 2'b01;
      12'h217: color = 2'b01;
      12'h218: color = 2'b01;
      12'h219: color = 2'b01;
      12'h21a: color = 2'b01;
      12'h21b: color = 2'b10;
      12'h21c: color = 2'b10;
      12'h21d: color = 2'b10;
      12'h21e: color = 2'b01;
      12'h21f: color = 2'b01;
      12'h220: color = 2'b10;
      12'h221: color = 2'b10;
      12'h222: color = 2'b10;
      12'h223: color = 2'b10;
      12'h224: color = 2'b10;
      12'h225: color = 2'b10;
      12'h226: color = 2'b10;
      12'h227: color = 2'b10;
      12'h228: color = 2'b10;
      12'h229: color = 2'b10;
      12'h22a: color = 2'b10;
      12'h22b: color = 2'b00;
      12'h22c: color = 2'b00;
      12'h22d: color = 2'b00;
      12'h22e: color = 2'b11;
      12'h22f: color = 2'b11;
      12'h230: color = 2'b11;
      12'h231: color = 2'b11;
      12'h232: color = 2'b11;
      12'h233: color = 2'b11;
      12'h234: color = 2'b11;
      12'h235: color = 2'b11;
      12'h236: color = 2'b11;
      12'h237: color = 2'b11;
      12'h238: color = 2'b11;
      12'h239: color = 2'b11;
      12'h23a: color = 2'b11;
      12'h23b: color = 2'b11;
      12'h23c: color = 2'b11;
      12'h23d: color = 2'b11;
      12'h23e: color = 2'b11;
      12'h23f: color = 2'b11;
      12'h240: color = 2'b11;
      12'h241: color = 2'b11;
      12'h242: color = 2'b11;
      12'h243: color = 2'b11;
      12'h244: color = 2'b11;
      12'h245: color = 2'b11;
      12'h246: color = 2'b11;
      12'h247: color = 2'b11;
      12'h248: color = 2'b11;
      12'h249: color = 2'b11;
      12'h24a: color = 2'b11;
      12'h24b: color = 2'b11;
      12'h24c: color = 2'b11;
      12'h24d: color = 2'b11;
      12'h24e: color = 2'b00;
      12'h24f: color = 2'b00;
      12'h250: color = 2'b01;
      12'h251: color = 2'b01;
      12'h252: color = 2'b01;
      12'h253: color = 2'b01;
      12'h254: color = 2'b01;
      12'h255: color = 2'b01;
      12'h256: color = 2'b01;
      12'h257: color = 2'b01;
      12'h258: color = 2'b01;
      12'h259: color = 2'b01;
      12'h25a: color = 2'b01;
      12'h25b: color = 2'b01;
      12'h25c: color = 2'b01;
      12'h25d: color = 2'b01;
      12'h25e: color = 2'b10;
      12'h25f: color = 2'b10;
      12'h260: color = 2'b01;
      12'h261: color = 2'b01;
      12'h262: color = 2'b10;
      12'h263: color = 2'b10;
      12'h264: color = 2'b10;
      12'h265: color = 2'b10;
      12'h266: color = 2'b10;
      12'h267: color = 2'b10;
      12'h268: color = 2'b10;
      12'h269: color = 2'b10;
      12'h26a: color = 2'b10;
      12'h26b: color = 2'b10;
      12'h26c: color = 2'b10;
      12'h26d: color = 2'b10;
      12'h26e: color = 2'b01;
      12'h26f: color = 2'b01;
      12'h270: color = 2'b11;
      12'h271: color = 2'b11;
      12'h272: color = 2'b11;
      12'h273: color = 2'b11;
      12'h274: color = 2'b11;
      12'h275: color = 2'b11;
      12'h276: color = 2'b11;
      12'h277: color = 2'b11;
      12'h278: color = 2'b11;
      12'h279: color = 2'b11;
      12'h27a: color = 2'b11;
      12'h27b: color = 2'b11;
      12'h27c: color = 2'b11;
      12'h27d: color = 2'b11;
      12'h27e: color = 2'b11;
      12'h27f: color = 2'b11;
      12'h280: color = 2'b11;
      12'h281: color = 2'b11;
      12'h282: color = 2'b11;
      12'h283: color = 2'b11;
      12'h284: color = 2'b11;
      12'h285: color = 2'b11;
      12'h286: color = 2'b11;
      12'h287: color = 2'b11;
      12'h288: color = 2'b11;
      12'h289: color = 2'b11;
      12'h28a: color = 2'b11;
      12'h28b: color = 2'b11;
      12'h28c: color = 2'b11;
      12'h28d: color = 2'b11;
      12'h28e: color = 2'b00;
      12'h28f: color = 2'b00;
      12'h290: color = 2'b01;
      12'h291: color = 2'b01;
      12'h292: color = 2'b01;
      12'h293: color = 2'b01;
      12'h294: color = 2'b01;
      12'h295: color = 2'b01;
      12'h296: color = 2'b01;
      12'h297: color = 2'b01;
      12'h298: color = 2'b01;
      12'h299: color = 2'b01;
      12'h29a: color = 2'b01;
      12'h29b: color = 2'b01;
      12'h29c: color = 2'b01;
      12'h29d: color = 2'b01;
      12'h29e: color = 2'b10;
      12'h29f: color = 2'b10;
      12'h2a0: color = 2'b01;
      12'h2a1: color = 2'b01;
      12'h2a2: color = 2'b10;
      12'h2a3: color = 2'b10;
      12'h2a4: color = 2'b10;
      12'h2a5: color = 2'b10;
      12'h2a6: color = 2'b10;
      12'h2a7: color = 2'b10;
      12'h2a8: color = 2'b10;
      12'h2a9: color = 2'b10;
      12'h2aa: color = 2'b10;
      12'h2ab: color = 2'b10;
      12'h2ac: color = 2'b10;
      12'h2ad: color = 2'b10;
      12'h2ae: color = 2'b01;
      12'h2af: color = 2'b01;
      12'h2b0: color = 2'b11;
      12'h2b1: color = 2'b11;
      12'h2b2: color = 2'b11;
      12'h2b3: color = 2'b11;
      12'h2b4: color = 2'b11;
      12'h2b5: color = 2'b11;
      12'h2b6: color = 2'b11;
      12'h2b7: color = 2'b11;
      12'h2b8: color = 2'b11;
      12'h2b9: color = 2'b11;
      12'h2ba: color = 2'b11;
      12'h2bb: color = 2'b11;
      12'h2bc: color = 2'b11;
      12'h2bd: color = 2'b11;
      12'h2be: color = 2'b11;
      12'h2bf: color = 2'b11;
      12'h2c0: color = 2'b11;
      12'h2c1: color = 2'b11;
      12'h2c2: color = 2'b11;
      12'h2c3: color = 2'b11;
      12'h2c4: color = 2'b11;
      12'h2c5: color = 2'b11;
      12'h2c6: color = 2'b11;
      12'h2c7: color = 2'b11;
      12'h2c8: color = 2'b11;
      12'h2c9: color = 2'b11;
      12'h2ca: color = 2'b11;
      12'h2cb: color = 2'b00;
      12'h2cc: color = 2'b00;
      12'h2cd: color = 2'b00;
      12'h2ce: color = 2'b01;
      12'h2cf: color = 2'b01;
      12'h2d0: color = 2'b01;
      12'h2d1: color = 2'b01;
      12'h2d2: color = 2'b01;
      12'h2d3: color = 2'b01;
      12'h2d4: color = 2'b01;
      12'h2d5: color = 2'b01;
      12'h2d6: color = 2'b01;
      12'h2d7: color = 2'b01;
      12'h2d8: color = 2'b01;
      12'h2d9: color = 2'b01;
      12'h2da: color = 2'b01;
      12'h2db: color = 2'b01;
      12'h2dc: color = 2'b01;
      12'h2dd: color = 2'b01;
      12'h2de: color = 2'b01;
      12'h2df: color = 2'b01;
      12'h2e0: color = 2'b10;
      12'h2e1: color = 2'b10;
      12'h2e2: color = 2'b01;
      12'h2e3: color = 2'b01;
      12'h2e4: color = 2'b01;
      12'h2e5: color = 2'b10;
      12'h2e6: color = 2'b10;
      12'h2e7: color = 2'b10;
      12'h2e8: color = 2'b10;
      12'h2e9: color = 2'b10;
      12'h2ea: color = 2'b10;
      12'h2eb: color = 2'b10;
      12'h2ec: color = 2'b10;
      12'h2ed: color = 2'b10;
      12'h2ee: color = 2'b00;
      12'h2ef: color = 2'b00;
      12'h2f0: color = 2'b11;
      12'h2f1: color = 2'b11;
      12'h2f2: color = 2'b11;
      12'h2f3: color = 2'b11;
      12'h2f4: color = 2'b11;
      12'h2f5: color = 2'b11;
      12'h2f6: color = 2'b11;
      12'h2f7: color = 2'b11;
      12'h2f8: color = 2'b11;
      12'h2f9: color = 2'b11;
      12'h2fa: color = 2'b11;
      12'h2fb: color = 2'b11;
      12'h2fc: color = 2'b11;
      12'h2fd: color = 2'b11;
      12'h2fe: color = 2'b11;
      12'h2ff: color = 2'b11;
      12'h300: color = 2'b11;
      12'h301: color = 2'b11;
      12'h302: color = 2'b11;
      12'h303: color = 2'b11;
      12'h304: color = 2'b11;
      12'h305: color = 2'b11;
      12'h306: color = 2'b11;
      12'h307: color = 2'b11;
      12'h308: color = 2'b11;
      12'h309: color = 2'b11;
      12'h30a: color = 2'b11;
      12'h30b: color = 2'b00;
      12'h30c: color = 2'b00;
      12'h30d: color = 2'b00;
      12'h30e: color = 2'b01;
      12'h30f: color = 2'b01;
      12'h310: color = 2'b01;
      12'h311: color = 2'b01;
      12'h312: color = 2'b01;
      12'h313: color = 2'b01;
      12'h314: color = 2'b01;
      12'h315: color = 2'b01;
      12'h316: color = 2'b01;
      12'h317: color = 2'b01;
      12'h318: color = 2'b01;
      12'h319: color = 2'b01;
      12'h31a: color = 2'b01;
      12'h31b: color = 2'b01;
      12'h31c: color = 2'b01;
      12'h31d: color = 2'b01;
      12'h31e: color = 2'b01;
      12'h31f: color = 2'b01;
      12'h320: color = 2'b10;
      12'h321: color = 2'b10;
      12'h322: color = 2'b01;
      12'h323: color = 2'b01;
      12'h324: color = 2'b01;
      12'h325: color = 2'b10;
      12'h326: color = 2'b10;
      12'h327: color = 2'b10;
      12'h328: color = 2'b10;
      12'h329: color = 2'b10;
      12'h32a: color = 2'b10;
      12'h32b: color = 2'b10;
      12'h32c: color = 2'b10;
      12'h32d: color = 2'b10;
      12'h32e: color = 2'b00;
      12'h32f: color = 2'b00;
      12'h330: color = 2'b11;
      12'h331: color = 2'b11;
      12'h332: color = 2'b11;
      12'h333: color = 2'b11;
      12'h334: color = 2'b11;
      12'h335: color = 2'b11;
      12'h336: color = 2'b11;
      12'h337: color = 2'b11;
      12'h338: color = 2'b11;
      12'h339: color = 2'b11;
      12'h33a: color = 2'b11;
      12'h33b: color = 2'b11;
      12'h33c: color = 2'b11;
      12'h33d: color = 2'b11;
      12'h33e: color = 2'b11;
      12'h33f: color = 2'b11;
      12'h340: color = 2'b11;
      12'h341: color = 2'b11;
      12'h342: color = 2'b11;
      12'h343: color = 2'b11;
      12'h344: color = 2'b11;
      12'h345: color = 2'b11;
      12'h346: color = 2'b11;
      12'h347: color = 2'b11;
      12'h348: color = 2'b11;
      12'h349: color = 2'b11;
      12'h34a: color = 2'b11;
      12'h34b: color = 2'b00;
      12'h34c: color = 2'b00;
      12'h34d: color = 2'b00;
      12'h34e: color = 2'b01;
      12'h34f: color = 2'b01;
      12'h350: color = 2'b01;
      12'h351: color = 2'b01;
      12'h352: color = 2'b01;
      12'h353: color = 2'b01;
      12'h354: color = 2'b01;
      12'h355: color = 2'b01;
      12'h356: color = 2'b01;
      12'h357: color = 2'b01;
      12'h358: color = 2'b01;
      12'h359: color = 2'b01;
      12'h35a: color = 2'b01;
      12'h35b: color = 2'b01;
      12'h35c: color = 2'b01;
      12'h35d: color = 2'b01;
      12'h35e: color = 2'b10;
      12'h35f: color = 2'b10;
      12'h360: color = 2'b01;
      12'h361: color = 2'b01;
      12'h362: color = 2'b10;
      12'h363: color = 2'b10;
      12'h364: color = 2'b10;
      12'h365: color = 2'b01;
      12'h366: color = 2'b01;
      12'h367: color = 2'b10;
      12'h368: color = 2'b10;
      12'h369: color = 2'b10;
      12'h36a: color = 2'b10;
      12'h36b: color = 2'b10;
      12'h36c: color = 2'b10;
      12'h36d: color = 2'b10;
      12'h36e: color = 2'b00;
      12'h36f: color = 2'b00;
      12'h370: color = 2'b00;
      12'h371: color = 2'b00;
      12'h372: color = 2'b00;
      12'h373: color = 2'b00;
      12'h374: color = 2'b00;
      12'h375: color = 2'b11;
      12'h376: color = 2'b11;
      12'h377: color = 2'b11;
      12'h378: color = 2'b11;
      12'h379: color = 2'b11;
      12'h37a: color = 2'b11;
      12'h37b: color = 2'b11;
      12'h37c: color = 2'b11;
      12'h37d: color = 2'b11;
      12'h37e: color = 2'b11;
      12'h37f: color = 2'b11;
      12'h380: color = 2'b11;
      12'h381: color = 2'b11;
      12'h382: color = 2'b11;
      12'h383: color = 2'b11;
      12'h384: color = 2'b11;
      12'h385: color = 2'b11;
      12'h386: color = 2'b11;
      12'h387: color = 2'b11;
      12'h388: color = 2'b11;
      12'h389: color = 2'b11;
      12'h38a: color = 2'b11;
      12'h38b: color = 2'b00;
      12'h38c: color = 2'b00;
      12'h38d: color = 2'b00;
      12'h38e: color = 2'b01;
      12'h38f: color = 2'b01;
      12'h390: color = 2'b01;
      12'h391: color = 2'b01;
      12'h392: color = 2'b01;
      12'h393: color = 2'b01;
      12'h394: color = 2'b01;
      12'h395: color = 2'b01;
      12'h396: color = 2'b01;
      12'h397: color = 2'b01;
      12'h398: color = 2'b01;
      12'h399: color = 2'b01;
      12'h39a: color = 2'b01;
      12'h39b: color = 2'b01;
      12'h39c: color = 2'b01;
      12'h39d: color = 2'b01;
      12'h39e: color = 2'b10;
      12'h39f: color = 2'b10;
      12'h3a0: color = 2'b01;
      12'h3a1: color = 2'b01;
      12'h3a2: color = 2'b10;
      12'h3a3: color = 2'b10;
      12'h3a4: color = 2'b10;
      12'h3a5: color = 2'b01;
      12'h3a6: color = 2'b01;
      12'h3a7: color = 2'b10;
      12'h3a8: color = 2'b10;
      12'h3a9: color = 2'b10;
      12'h3aa: color = 2'b10;
      12'h3ab: color = 2'b10;
      12'h3ac: color = 2'b10;
      12'h3ad: color = 2'b10;
      12'h3ae: color = 2'b00;
      12'h3af: color = 2'b00;
      12'h3b0: color = 2'b00;
      12'h3b1: color = 2'b00;
      12'h3b2: color = 2'b00;
      12'h3b3: color = 2'b00;
      12'h3b4: color = 2'b00;
      12'h3b5: color = 2'b11;
      12'h3b6: color = 2'b11;
      12'h3b7: color = 2'b11;
      12'h3b8: color = 2'b11;
      12'h3b9: color = 2'b11;
      12'h3ba: color = 2'b11;
      12'h3bb: color = 2'b11;
      12'h3bc: color = 2'b11;
      12'h3bd: color = 2'b11;
      12'h3be: color = 2'b11;
      12'h3bf: color = 2'b11;
      12'h3c0: color = 2'b11;
      12'h3c1: color = 2'b11;
      12'h3c2: color = 2'b11;
      12'h3c3: color = 2'b11;
      12'h3c4: color = 2'b11;
      12'h3c5: color = 2'b11;
      12'h3c6: color = 2'b11;
      12'h3c7: color = 2'b11;
      12'h3c8: color = 2'b11;
      12'h3c9: color = 2'b11;
      12'h3ca: color = 2'b11;
      12'h3cb: color = 2'b00;
      12'h3cc: color = 2'b00;
      12'h3cd: color = 2'b00;
      12'h3ce: color = 2'b01;
      12'h3cf: color = 2'b01;
      12'h3d0: color = 2'b01;
      12'h3d1: color = 2'b01;
      12'h3d2: color = 2'b01;
      12'h3d3: color = 2'b01;
      12'h3d4: color = 2'b01;
      12'h3d5: color = 2'b01;
      12'h3d6: color = 2'b01;
      12'h3d7: color = 2'b01;
      12'h3d8: color = 2'b01;
      12'h3d9: color = 2'b01;
      12'h3da: color = 2'b01;
      12'h3db: color = 2'b01;
      12'h3dc: color = 2'b01;
      12'h3dd: color = 2'b01;
      12'h3de: color = 2'b10;
      12'h3df: color = 2'b10;
      12'h3e0: color = 2'b01;
      12'h3e1: color = 2'b01;
      12'h3e2: color = 2'b10;
      12'h3e3: color = 2'b10;
      12'h3e4: color = 2'b10;
      12'h3e5: color = 2'b01;
      12'h3e6: color = 2'b01;
      12'h3e7: color = 2'b10;
      12'h3e8: color = 2'b10;
      12'h3e9: color = 2'b10;
      12'h3ea: color = 2'b10;
      12'h3eb: color = 2'b10;
      12'h3ec: color = 2'b10;
      12'h3ed: color = 2'b10;
      12'h3ee: color = 2'b00;
      12'h3ef: color = 2'b00;
      12'h3f0: color = 2'b00;
      12'h3f1: color = 2'b00;
      12'h3f2: color = 2'b00;
      12'h3f3: color = 2'b00;
      12'h3f4: color = 2'b00;
      12'h3f5: color = 2'b11;
      12'h3f6: color = 2'b11;
      12'h3f7: color = 2'b11;
      12'h3f8: color = 2'b11;
      12'h3f9: color = 2'b11;
      12'h3fa: color = 2'b11;
      12'h3fb: color = 2'b11;
      12'h3fc: color = 2'b11;
      12'h3fd: color = 2'b11;
      12'h3fe: color = 2'b11;
      12'h3ff: color = 2'b11;
      12'h400: color = 2'b11;
      12'h401: color = 2'b11;
      12'h402: color = 2'b11;
      12'h403: color = 2'b11;
      12'h404: color = 2'b11;
      12'h405: color = 2'b11;
      12'h406: color = 2'b11;
      12'h407: color = 2'b11;
      12'h408: color = 2'b11;
      12'h409: color = 2'b11;
      12'h40a: color = 2'b11;
      12'h40b: color = 2'b00;
      12'h40c: color = 2'b00;
      12'h40d: color = 2'b00;
      12'h40e: color = 2'b01;
      12'h40f: color = 2'b01;
      12'h410: color = 2'b01;
      12'h411: color = 2'b01;
      12'h412: color = 2'b01;
      12'h413: color = 2'b01;
      12'h414: color = 2'b01;
      12'h415: color = 2'b01;
      12'h416: color = 2'b01;
      12'h417: color = 2'b01;
      12'h418: color = 2'b01;
      12'h419: color = 2'b01;
      12'h41a: color = 2'b01;
      12'h41b: color = 2'b01;
      12'h41c: color = 2'b01;
      12'h41d: color = 2'b01;
      12'h41e: color = 2'b01;
      12'h41f: color = 2'b01;
      12'h420: color = 2'b01;
      12'h421: color = 2'b01;
      12'h422: color = 2'b01;
      12'h423: color = 2'b01;
      12'h424: color = 2'b01;
      12'h425: color = 2'b01;
      12'h426: color = 2'b01;
      12'h427: color = 2'b01;
      12'h428: color = 2'b01;
      12'h429: color = 2'b01;
      12'h42a: color = 2'b01;
      12'h42b: color = 2'b11;
      12'h42c: color = 2'b11;
      12'h42d: color = 2'b11;
      12'h42e: color = 2'b11;
      12'h42f: color = 2'b11;
      12'h430: color = 2'b11;
      12'h431: color = 2'b11;
      12'h432: color = 2'b11;
      12'h433: color = 2'b11;
      12'h434: color = 2'b11;
      12'h435: color = 2'b00;
      12'h436: color = 2'b00;
      12'h437: color = 2'b11;
      12'h438: color = 2'b11;
      12'h439: color = 2'b11;
      12'h43a: color = 2'b11;
      12'h43b: color = 2'b11;
      12'h43c: color = 2'b11;
      12'h43d: color = 2'b11;
      12'h43e: color = 2'b11;
      12'h43f: color = 2'b11;
      12'h440: color = 2'b11;
      12'h441: color = 2'b11;
      12'h442: color = 2'b11;
      12'h443: color = 2'b11;
      12'h444: color = 2'b11;
      12'h445: color = 2'b11;
      12'h446: color = 2'b11;
      12'h447: color = 2'b11;
      12'h448: color = 2'b11;
      12'h449: color = 2'b11;
      12'h44a: color = 2'b11;
      12'h44b: color = 2'b00;
      12'h44c: color = 2'b00;
      12'h44d: color = 2'b00;
      12'h44e: color = 2'b01;
      12'h44f: color = 2'b01;
      12'h450: color = 2'b01;
      12'h451: color = 2'b01;
      12'h452: color = 2'b01;
      12'h453: color = 2'b01;
      12'h454: color = 2'b01;
      12'h455: color = 2'b01;
      12'h456: color = 2'b01;
      12'h457: color = 2'b01;
      12'h458: color = 2'b01;
      12'h459: color = 2'b01;
      12'h45a: color = 2'b01;
      12'h45b: color = 2'b01;
      12'h45c: color = 2'b01;
      12'h45d: color = 2'b01;
      12'h45e: color = 2'b01;
      12'h45f: color = 2'b01;
      12'h460: color = 2'b01;
      12'h461: color = 2'b01;
      12'h462: color = 2'b01;
      12'h463: color = 2'b01;
      12'h464: color = 2'b01;
      12'h465: color = 2'b01;
      12'h466: color = 2'b01;
      12'h467: color = 2'b01;
      12'h468: color = 2'b01;
      12'h469: color = 2'b01;
      12'h46a: color = 2'b01;
      12'h46b: color = 2'b11;
      12'h46c: color = 2'b11;
      12'h46d: color = 2'b11;
      12'h46e: color = 2'b11;
      12'h46f: color = 2'b11;
      12'h470: color = 2'b11;
      12'h471: color = 2'b11;
      12'h472: color = 2'b11;
      12'h473: color = 2'b11;
      12'h474: color = 2'b11;
      12'h475: color = 2'b00;
      12'h476: color = 2'b00;
      12'h477: color = 2'b11;
      12'h478: color = 2'b11;
      12'h479: color = 2'b11;
      12'h47a: color = 2'b11;
      12'h47b: color = 2'b11;
      12'h47c: color = 2'b11;
      12'h47d: color = 2'b11;
      12'h47e: color = 2'b11;
      12'h47f: color = 2'b11;
      12'h480: color = 2'b11;
      12'h481: color = 2'b11;
      12'h482: color = 2'b11;
      12'h483: color = 2'b11;
      12'h484: color = 2'b11;
      12'h485: color = 2'b11;
      12'h486: color = 2'b11;
      12'h487: color = 2'b11;
      12'h488: color = 2'b11;
      12'h489: color = 2'b11;
      12'h48a: color = 2'b11;
      12'h48b: color = 2'b11;
      12'h48c: color = 2'b11;
      12'h48d: color = 2'b11;
      12'h48e: color = 2'b01;
      12'h48f: color = 2'b01;
      12'h490: color = 2'b01;
      12'h491: color = 2'b01;
      12'h492: color = 2'b00;
      12'h493: color = 2'b00;
      12'h494: color = 2'b00;
      12'h495: color = 2'b00;
      12'h496: color = 2'b00;
      12'h497: color = 2'b00;
      12'h498: color = 2'b00;
      12'h499: color = 2'b01;
      12'h49a: color = 2'b01;
      12'h49b: color = 2'b01;
      12'h49c: color = 2'b01;
      12'h49d: color = 2'b01;
      12'h49e: color = 2'b01;
      12'h49f: color = 2'b01;
      12'h4a0: color = 2'b01;
      12'h4a1: color = 2'b01;
      12'h4a2: color = 2'b01;
      12'h4a3: color = 2'b01;
      12'h4a4: color = 2'b01;
      12'h4a5: color = 2'b01;
      12'h4a6: color = 2'b01;
      12'h4a7: color = 2'b11;
      12'h4a8: color = 2'b11;
      12'h4a9: color = 2'b11;
      12'h4aa: color = 2'b11;
      12'h4ab: color = 2'b11;
      12'h4ac: color = 2'b11;
      12'h4ad: color = 2'b11;
      12'h4ae: color = 2'b11;
      12'h4af: color = 2'b11;
      12'h4b0: color = 2'b00;
      12'h4b1: color = 2'b00;
      12'h4b2: color = 2'b00;
      12'h4b3: color = 2'b00;
      12'h4b4: color = 2'b00;
      12'h4b5: color = 2'b11;
      12'h4b6: color = 2'b11;
      12'h4b7: color = 2'b11;
      12'h4b8: color = 2'b11;
      12'h4b9: color = 2'b11;
      12'h4ba: color = 2'b11;
      12'h4bb: color = 2'b11;
      12'h4bc: color = 2'b11;
      12'h4bd: color = 2'b11;
      12'h4be: color = 2'b11;
      12'h4bf: color = 2'b11;
      12'h4c0: color = 2'b11;
      12'h4c1: color = 2'b11;
      12'h4c2: color = 2'b11;
      12'h4c3: color = 2'b11;
      12'h4c4: color = 2'b11;
      12'h4c5: color = 2'b11;
      12'h4c6: color = 2'b11;
      12'h4c7: color = 2'b11;
      12'h4c8: color = 2'b11;
      12'h4c9: color = 2'b11;
      12'h4ca: color = 2'b11;
      12'h4cb: color = 2'b11;
      12'h4cc: color = 2'b11;
      12'h4cd: color = 2'b11;
      12'h4ce: color = 2'b01;
      12'h4cf: color = 2'b01;
      12'h4d0: color = 2'b01;
      12'h4d1: color = 2'b01;
      12'h4d2: color = 2'b00;
      12'h4d3: color = 2'b00;
      12'h4d4: color = 2'b00;
      12'h4d5: color = 2'b00;
      12'h4d6: color = 2'b00;
      12'h4d7: color = 2'b00;
      12'h4d8: color = 2'b00;
      12'h4d9: color = 2'b01;
      12'h4da: color = 2'b01;
      12'h4db: color = 2'b01;
      12'h4dc: color = 2'b01;
      12'h4dd: color = 2'b01;
      12'h4de: color = 2'b01;
      12'h4df: color = 2'b01;
      12'h4e0: color = 2'b01;
      12'h4e1: color = 2'b01;
      12'h4e2: color = 2'b01;
      12'h4e3: color = 2'b01;
      12'h4e4: color = 2'b01;
      12'h4e5: color = 2'b01;
      12'h4e6: color = 2'b01;
      12'h4e7: color = 2'b11;
      12'h4e8: color = 2'b11;
      12'h4e9: color = 2'b11;
      12'h4ea: color = 2'b11;
      12'h4eb: color = 2'b11;
      12'h4ec: color = 2'b11;
      12'h4ed: color = 2'b11;
      12'h4ee: color = 2'b11;
      12'h4ef: color = 2'b11;
      12'h4f0: color = 2'b00;
      12'h4f1: color = 2'b00;
      12'h4f2: color = 2'b00;
      12'h4f3: color = 2'b00;
      12'h4f4: color = 2'b00;
      12'h4f5: color = 2'b11;
      12'h4f6: color = 2'b11;
      12'h4f7: color = 2'b11;
      12'h4f8: color = 2'b11;
      12'h4f9: color = 2'b11;
      12'h4fa: color = 2'b11;
      12'h4fb: color = 2'b11;
      12'h4fc: color = 2'b11;
      12'h4fd: color = 2'b11;
      12'h4fe: color = 2'b11;
      12'h4ff: color = 2'b11;
      12'h500: color = 2'b11;
      12'h501: color = 2'b11;
      12'h502: color = 2'b11;
      12'h503: color = 2'b11;
      12'h504: color = 2'b11;
      12'h505: color = 2'b11;
      12'h506: color = 2'b11;
      12'h507: color = 2'b11;
      12'h508: color = 2'b11;
      12'h509: color = 2'b11;
      12'h50a: color = 2'b11;
      12'h50b: color = 2'b11;
      12'h50c: color = 2'b11;
      12'h50d: color = 2'b11;
      12'h50e: color = 2'b00;
      12'h50f: color = 2'b00;
      12'h510: color = 2'b01;
      12'h511: color = 2'b01;
      12'h512: color = 2'b01;
      12'h513: color = 2'b01;
      12'h514: color = 2'b01;
      12'h515: color = 2'b01;
      12'h516: color = 2'b01;
      12'h517: color = 2'b01;
      12'h518: color = 2'b01;
      12'h519: color = 2'b01;
      12'h51a: color = 2'b01;
      12'h51b: color = 2'b01;
      12'h51c: color = 2'b01;
      12'h51d: color = 2'b01;
      12'h51e: color = 2'b01;
      12'h51f: color = 2'b01;
      12'h520: color = 2'b00;
      12'h521: color = 2'b00;
      12'h522: color = 2'b00;
      12'h523: color = 2'b00;
      12'h524: color = 2'b00;
      12'h525: color = 2'b00;
      12'h526: color = 2'b00;
      12'h527: color = 2'b01;
      12'h528: color = 2'b01;
      12'h529: color = 2'b01;
      12'h52a: color = 2'b01;
      12'h52b: color = 2'b00;
      12'h52c: color = 2'b00;
      12'h52d: color = 2'b00;
      12'h52e: color = 2'b00;
      12'h52f: color = 2'b00;
      12'h530: color = 2'b11;
      12'h531: color = 2'b11;
      12'h532: color = 2'b11;
      12'h533: color = 2'b11;
      12'h534: color = 2'b11;
      12'h535: color = 2'b11;
      12'h536: color = 2'b11;
      12'h537: color = 2'b11;
      12'h538: color = 2'b11;
      12'h539: color = 2'b11;
      12'h53a: color = 2'b11;
      12'h53b: color = 2'b11;
      12'h53c: color = 2'b11;
      12'h53d: color = 2'b11;
      12'h53e: color = 2'b11;
      12'h53f: color = 2'b11;
      12'h540: color = 2'b11;
      12'h541: color = 2'b11;
      12'h542: color = 2'b11;
      12'h543: color = 2'b11;
      12'h544: color = 2'b11;
      12'h545: color = 2'b11;
      12'h546: color = 2'b11;
      12'h547: color = 2'b11;
      12'h548: color = 2'b11;
      12'h549: color = 2'b11;
      12'h54a: color = 2'b11;
      12'h54b: color = 2'b11;
      12'h54c: color = 2'b11;
      12'h54d: color = 2'b11;
      12'h54e: color = 2'b00;
      12'h54f: color = 2'b00;
      12'h550: color = 2'b01;
      12'h551: color = 2'b01;
      12'h552: color = 2'b01;
      12'h553: color = 2'b01;
      12'h554: color = 2'b01;
      12'h555: color = 2'b01;
      12'h556: color = 2'b01;
      12'h557: color = 2'b01;
      12'h558: color = 2'b01;
      12'h559: color = 2'b01;
      12'h55a: color = 2'b01;
      12'h55b: color = 2'b01;
      12'h55c: color = 2'b01;
      12'h55d: color = 2'b01;
      12'h55e: color = 2'b01;
      12'h55f: color = 2'b01;
      12'h560: color = 2'b00;
      12'h561: color = 2'b00;
      12'h562: color = 2'b00;
      12'h563: color = 2'b00;
      12'h564: color = 2'b00;
      12'h565: color = 2'b00;
      12'h566: color = 2'b00;
      12'h567: color = 2'b01;
      12'h568: color = 2'b01;
      12'h569: color = 2'b01;
      12'h56a: color = 2'b01;
      12'h56b: color = 2'b00;
      12'h56c: color = 2'b00;
      12'h56d: color = 2'b00;
      12'h56e: color = 2'b00;
      12'h56f: color = 2'b00;
      12'h570: color = 2'b11;
      12'h571: color = 2'b11;
      12'h572: color = 2'b11;
      12'h573: color = 2'b11;
      12'h574: color = 2'b11;
      12'h575: color = 2'b11;
      12'h576: color = 2'b11;
      12'h577: color = 2'b11;
      12'h578: color = 2'b11;
      12'h579: color = 2'b11;
      12'h57a: color = 2'b11;
      12'h57b: color = 2'b11;
      12'h57c: color = 2'b11;
      12'h57d: color = 2'b11;
      12'h57e: color = 2'b11;
      12'h57f: color = 2'b11;
      12'h580: color = 2'b11;
      12'h581: color = 2'b11;
      12'h582: color = 2'b11;
      12'h583: color = 2'b11;
      12'h584: color = 2'b11;
      12'h585: color = 2'b11;
      12'h586: color = 2'b11;
      12'h587: color = 2'b11;
      12'h588: color = 2'b11;
      12'h589: color = 2'b11;
      12'h58a: color = 2'b11;
      12'h58b: color = 2'b11;
      12'h58c: color = 2'b11;
      12'h58d: color = 2'b11;
      12'h58e: color = 2'b00;
      12'h58f: color = 2'b00;
      12'h590: color = 2'b00;
      12'h591: color = 2'b00;
      12'h592: color = 2'b00;
      12'h593: color = 2'b00;
      12'h594: color = 2'b00;
      12'h595: color = 2'b00;
      12'h596: color = 2'b00;
      12'h597: color = 2'b00;
      12'h598: color = 2'b00;
      12'h599: color = 2'b00;
      12'h59a: color = 2'b00;
      12'h59b: color = 2'b00;
      12'h59c: color = 2'b00;
      12'h59d: color = 2'b00;
      12'h59e: color = 2'b00;
      12'h59f: color = 2'b00;
      12'h5a0: color = 2'b00;
      12'h5a1: color = 2'b00;
      12'h5a2: color = 2'b00;
      12'h5a3: color = 2'b00;
      12'h5a4: color = 2'b00;
      12'h5a5: color = 2'b11;
      12'h5a6: color = 2'b11;
      12'h5a7: color = 2'b00;
      12'h5a8: color = 2'b00;
      12'h5a9: color = 2'b10;
      12'h5aa: color = 2'b10;
      12'h5ab: color = 2'b00;
      12'h5ac: color = 2'b00;
      12'h5ad: color = 2'b00;
      12'h5ae: color = 2'b00;
      12'h5af: color = 2'b00;
      12'h5b0: color = 2'b11;
      12'h5b1: color = 2'b11;
      12'h5b2: color = 2'b11;
      12'h5b3: color = 2'b11;
      12'h5b4: color = 2'b11;
      12'h5b5: color = 2'b11;
      12'h5b6: color = 2'b11;
      12'h5b7: color = 2'b11;
      12'h5b8: color = 2'b11;
      12'h5b9: color = 2'b11;
      12'h5ba: color = 2'b11;
      12'h5bb: color = 2'b11;
      12'h5bc: color = 2'b11;
      12'h5bd: color = 2'b11;
      12'h5be: color = 2'b11;
      12'h5bf: color = 2'b11;
      12'h5c0: color = 2'b11;
      12'h5c1: color = 2'b11;
      12'h5c2: color = 2'b11;
      12'h5c3: color = 2'b11;
      12'h5c4: color = 2'b11;
      12'h5c5: color = 2'b11;
      12'h5c6: color = 2'b11;
      12'h5c7: color = 2'b11;
      12'h5c8: color = 2'b11;
      12'h5c9: color = 2'b11;
      12'h5ca: color = 2'b11;
      12'h5cb: color = 2'b11;
      12'h5cc: color = 2'b11;
      12'h5cd: color = 2'b11;
      12'h5ce: color = 2'b00;
      12'h5cf: color = 2'b00;
      12'h5d0: color = 2'b00;
      12'h5d1: color = 2'b00;
      12'h5d2: color = 2'b00;
      12'h5d3: color = 2'b00;
      12'h5d4: color = 2'b00;
      12'h5d5: color = 2'b00;
      12'h5d6: color = 2'b00;
      12'h5d7: color = 2'b00;
      12'h5d8: color = 2'b00;
      12'h5d9: color = 2'b00;
      12'h5da: color = 2'b00;
      12'h5db: color = 2'b00;
      12'h5dc: color = 2'b00;
      12'h5dd: color = 2'b00;
      12'h5de: color = 2'b00;
      12'h5df: color = 2'b00;
      12'h5e0: color = 2'b00;
      12'h5e1: color = 2'b00;
      12'h5e2: color = 2'b00;
      12'h5e3: color = 2'b00;
      12'h5e4: color = 2'b00;
      12'h5e5: color = 2'b11;
      12'h5e6: color = 2'b11;
      12'h5e7: color = 2'b00;
      12'h5e8: color = 2'b00;
      12'h5e9: color = 2'b10;
      12'h5ea: color = 2'b10;
      12'h5eb: color = 2'b00;
      12'h5ec: color = 2'b00;
      12'h5ed: color = 2'b00;
      12'h5ee: color = 2'b00;
      12'h5ef: color = 2'b00;
      12'h5f0: color = 2'b11;
      12'h5f1: color = 2'b11;
      12'h5f2: color = 2'b11;
      12'h5f3: color = 2'b11;
      12'h5f4: color = 2'b11;
      12'h5f5: color = 2'b11;
      12'h5f6: color = 2'b11;
      12'h5f7: color = 2'b11;
      12'h5f8: color = 2'b11;
      12'h5f9: color = 2'b11;
      12'h5fa: color = 2'b11;
      12'h5fb: color = 2'b11;
      12'h5fc: color = 2'b11;
      12'h5fd: color = 2'b11;
      12'h5fe: color = 2'b11;
      12'h5ff: color = 2'b11;
      12'h600: color = 2'b11;
      12'h601: color = 2'b11;
      12'h602: color = 2'b11;
      12'h603: color = 2'b11;
      12'h604: color = 2'b11;
      12'h605: color = 2'b11;
      12'h606: color = 2'b11;
      12'h607: color = 2'b11;
      12'h608: color = 2'b11;
      12'h609: color = 2'b11;
      12'h60a: color = 2'b11;
      12'h60b: color = 2'b11;
      12'h60c: color = 2'b11;
      12'h60d: color = 2'b11;
      12'h60e: color = 2'b00;
      12'h60f: color = 2'b00;
      12'h610: color = 2'b00;
      12'h611: color = 2'b00;
      12'h612: color = 2'b00;
      12'h613: color = 2'b00;
      12'h614: color = 2'b00;
      12'h615: color = 2'b00;
      12'h616: color = 2'b00;
      12'h617: color = 2'b00;
      12'h618: color = 2'b00;
      12'h619: color = 2'b00;
      12'h61a: color = 2'b00;
      12'h61b: color = 2'b00;
      12'h61c: color = 2'b00;
      12'h61d: color = 2'b00;
      12'h61e: color = 2'b00;
      12'h61f: color = 2'b00;
      12'h620: color = 2'b00;
      12'h621: color = 2'b00;
      12'h622: color = 2'b00;
      12'h623: color = 2'b00;
      12'h624: color = 2'b00;
      12'h625: color = 2'b11;
      12'h626: color = 2'b11;
      12'h627: color = 2'b00;
      12'h628: color = 2'b00;
      12'h629: color = 2'b10;
      12'h62a: color = 2'b10;
      12'h62b: color = 2'b00;
      12'h62c: color = 2'b00;
      12'h62d: color = 2'b00;
      12'h62e: color = 2'b00;
      12'h62f: color = 2'b00;
      12'h630: color = 2'b11;
      12'h631: color = 2'b11;
      12'h632: color = 2'b11;
      12'h633: color = 2'b11;
      12'h634: color = 2'b11;
      12'h635: color = 2'b11;
      12'h636: color = 2'b11;
      12'h637: color = 2'b11;
      12'h638: color = 2'b11;
      12'h639: color = 2'b11;
      12'h63a: color = 2'b11;
      12'h63b: color = 2'b11;
      12'h63c: color = 2'b11;
      12'h63d: color = 2'b11;
      12'h63e: color = 2'b11;
      12'h63f: color = 2'b11;
      12'h640: color = 2'b11;
      12'h641: color = 2'b11;
      12'h642: color = 2'b11;
      12'h643: color = 2'b11;
      12'h644: color = 2'b11;
      12'h645: color = 2'b11;
      12'h646: color = 2'b11;
      12'h647: color = 2'b11;
      12'h648: color = 2'b11;
      12'h649: color = 2'b11;
      12'h64a: color = 2'b11;
      12'h64b: color = 2'b11;
      12'h64c: color = 2'b11;
      12'h64d: color = 2'b11;
      12'h64e: color = 2'b00;
      12'h64f: color = 2'b00;
      12'h650: color = 2'b00;
      12'h651: color = 2'b00;
      12'h652: color = 2'b00;
      12'h653: color = 2'b00;
      12'h654: color = 2'b00;
      12'h655: color = 2'b00;
      12'h656: color = 2'b00;
      12'h657: color = 2'b00;
      12'h658: color = 2'b00;
      12'h659: color = 2'b00;
      12'h65a: color = 2'b00;
      12'h65b: color = 2'b00;
      12'h65c: color = 2'b00;
      12'h65d: color = 2'b00;
      12'h65e: color = 2'b00;
      12'h65f: color = 2'b00;
      12'h660: color = 2'b00;
      12'h661: color = 2'b00;
      12'h662: color = 2'b00;
      12'h663: color = 2'b00;
      12'h664: color = 2'b00;
      12'h665: color = 2'b10;
      12'h666: color = 2'b10;
      12'h667: color = 2'b00;
      12'h668: color = 2'b00;
      12'h669: color = 2'b11;
      12'h66a: color = 2'b11;
      12'h66b: color = 2'b00;
      12'h66c: color = 2'b00;
      12'h66d: color = 2'b00;
      12'h66e: color = 2'b11;
      12'h66f: color = 2'b11;
      12'h670: color = 2'b11;
      12'h671: color = 2'b11;
      12'h672: color = 2'b11;
      12'h673: color = 2'b11;
      12'h674: color = 2'b11;
      12'h675: color = 2'b11;
      12'h676: color = 2'b11;
      12'h677: color = 2'b11;
      12'h678: color = 2'b11;
      12'h679: color = 2'b11;
      12'h67a: color = 2'b11;
      12'h67b: color = 2'b11;
      12'h67c: color = 2'b11;
      12'h67d: color = 2'b11;
      12'h67e: color = 2'b11;
      12'h67f: color = 2'b11;
      12'h680: color = 2'b11;
      12'h681: color = 2'b11;
      12'h682: color = 2'b11;
      12'h683: color = 2'b11;
      12'h684: color = 2'b11;
      12'h685: color = 2'b11;
      12'h686: color = 2'b11;
      12'h687: color = 2'b11;
      12'h688: color = 2'b11;
      12'h689: color = 2'b11;
      12'h68a: color = 2'b11;
      12'h68b: color = 2'b11;
      12'h68c: color = 2'b11;
      12'h68d: color = 2'b11;
      12'h68e: color = 2'b00;
      12'h68f: color = 2'b00;
      12'h690: color = 2'b00;
      12'h691: color = 2'b00;
      12'h692: color = 2'b00;
      12'h693: color = 2'b00;
      12'h694: color = 2'b00;
      12'h695: color = 2'b00;
      12'h696: color = 2'b00;
      12'h697: color = 2'b00;
      12'h698: color = 2'b00;
      12'h699: color = 2'b00;
      12'h69a: color = 2'b00;
      12'h69b: color = 2'b00;
      12'h69c: color = 2'b00;
      12'h69d: color = 2'b00;
      12'h69e: color = 2'b00;
      12'h69f: color = 2'b00;
      12'h6a0: color = 2'b00;
      12'h6a1: color = 2'b00;
      12'h6a2: color = 2'b00;
      12'h6a3: color = 2'b00;
      12'h6a4: color = 2'b00;
      12'h6a5: color = 2'b10;
      12'h6a6: color = 2'b10;
      12'h6a7: color = 2'b00;
      12'h6a8: color = 2'b00;
      12'h6a9: color = 2'b11;
      12'h6aa: color = 2'b11;
      12'h6ab: color = 2'b00;
      12'h6ac: color = 2'b00;
      12'h6ad: color = 2'b00;
      12'h6ae: color = 2'b11;
      12'h6af: color = 2'b11;
      12'h6b0: color = 2'b11;
      12'h6b1: color = 2'b11;
      12'h6b2: color = 2'b11;
      12'h6b3: color = 2'b11;
      12'h6b4: color = 2'b11;
      12'h6b5: color = 2'b11;
      12'h6b6: color = 2'b11;
      12'h6b7: color = 2'b11;
      12'h6b8: color = 2'b11;
      12'h6b9: color = 2'b11;
      12'h6ba: color = 2'b11;
      12'h6bb: color = 2'b11;
      12'h6bc: color = 2'b11;
      12'h6bd: color = 2'b11;
      12'h6be: color = 2'b11;
      12'h6bf: color = 2'b11;
      12'h6c0: color = 2'b11;
      12'h6c1: color = 2'b11;
      12'h6c2: color = 2'b11;
      12'h6c3: color = 2'b11;
      12'h6c4: color = 2'b11;
      12'h6c5: color = 2'b11;
      12'h6c6: color = 2'b11;
      12'h6c7: color = 2'b11;
      12'h6c8: color = 2'b11;
      12'h6c9: color = 2'b11;
      12'h6ca: color = 2'b11;
      12'h6cb: color = 2'b11;
      12'h6cc: color = 2'b11;
      12'h6cd: color = 2'b11;
      12'h6ce: color = 2'b11;
      12'h6cf: color = 2'b11;
      12'h6d0: color = 2'b00;
      12'h6d1: color = 2'b00;
      12'h6d2: color = 2'b00;
      12'h6d3: color = 2'b00;
      12'h6d4: color = 2'b00;
      12'h6d5: color = 2'b00;
      12'h6d6: color = 2'b00;
      12'h6d7: color = 2'b00;
      12'h6d8: color = 2'b00;
      12'h6d9: color = 2'b00;
      12'h6da: color = 2'b00;
      12'h6db: color = 2'b00;
      12'h6dc: color = 2'b00;
      12'h6dd: color = 2'b00;
      12'h6de: color = 2'b00;
      12'h6df: color = 2'b00;
      12'h6e0: color = 2'b00;
      12'h6e1: color = 2'b00;
      12'h6e2: color = 2'b00;
      12'h6e3: color = 2'b00;
      12'h6e4: color = 2'b00;
      12'h6e5: color = 2'b10;
      12'h6e6: color = 2'b10;
      12'h6e7: color = 2'b00;
      12'h6e8: color = 2'b00;
      12'h6e9: color = 2'b11;
      12'h6ea: color = 2'b11;
      12'h6eb: color = 2'b11;
      12'h6ec: color = 2'b11;
      12'h6ed: color = 2'b11;
      12'h6ee: color = 2'b01;
      12'h6ef: color = 2'b01;
      12'h6f0: color = 2'b11;
      12'h6f1: color = 2'b11;
      12'h6f2: color = 2'b11;
      12'h6f3: color = 2'b11;
      12'h6f4: color = 2'b11;
      12'h6f5: color = 2'b11;
      12'h6f6: color = 2'b11;
      12'h6f7: color = 2'b11;
      12'h6f8: color = 2'b11;
      12'h6f9: color = 2'b11;
      12'h6fa: color = 2'b11;
      12'h6fb: color = 2'b11;
      12'h6fc: color = 2'b11;
      12'h6fd: color = 2'b11;
      12'h6fe: color = 2'b11;
      12'h6ff: color = 2'b11;
      12'h700: color = 2'b11;
      12'h701: color = 2'b11;
      12'h702: color = 2'b11;
      12'h703: color = 2'b11;
      12'h704: color = 2'b11;
      12'h705: color = 2'b11;
      12'h706: color = 2'b11;
      12'h707: color = 2'b11;
      12'h708: color = 2'b11;
      12'h709: color = 2'b11;
      12'h70a: color = 2'b11;
      12'h70b: color = 2'b11;
      12'h70c: color = 2'b11;
      12'h70d: color = 2'b11;
      12'h70e: color = 2'b11;
      12'h70f: color = 2'b11;
      12'h710: color = 2'b00;
      12'h711: color = 2'b00;
      12'h712: color = 2'b00;
      12'h713: color = 2'b00;
      12'h714: color = 2'b00;
      12'h715: color = 2'b00;
      12'h716: color = 2'b00;
      12'h717: color = 2'b00;
      12'h718: color = 2'b00;
      12'h719: color = 2'b00;
      12'h71a: color = 2'b00;
      12'h71b: color = 2'b00;
      12'h71c: color = 2'b00;
      12'h71d: color = 2'b00;
      12'h71e: color = 2'b00;
      12'h71f: color = 2'b00;
      12'h720: color = 2'b00;
      12'h721: color = 2'b00;
      12'h722: color = 2'b00;
      12'h723: color = 2'b00;
      12'h724: color = 2'b00;
      12'h725: color = 2'b10;
      12'h726: color = 2'b10;
      12'h727: color = 2'b00;
      12'h728: color = 2'b00;
      12'h729: color = 2'b11;
      12'h72a: color = 2'b11;
      12'h72b: color = 2'b11;
      12'h72c: color = 2'b11;
      12'h72d: color = 2'b11;
      12'h72e: color = 2'b01;
      12'h72f: color = 2'b01;
      12'h730: color = 2'b11;
      12'h731: color = 2'b11;
      12'h732: color = 2'b11;
      12'h733: color = 2'b11;
      12'h734: color = 2'b11;
      12'h735: color = 2'b11;
      12'h736: color = 2'b11;
      12'h737: color = 2'b11;
      12'h738: color = 2'b11;
      12'h739: color = 2'b11;
      12'h73a: color = 2'b11;
      12'h73b: color = 2'b11;
      12'h73c: color = 2'b11;
      12'h73d: color = 2'b11;
      12'h73e: color = 2'b11;
      12'h73f: color = 2'b11;
      12'h740: color = 2'b11;
      12'h741: color = 2'b11;
      12'h742: color = 2'b11;
      12'h743: color = 2'b11;
      12'h744: color = 2'b11;
      12'h745: color = 2'b11;
      12'h746: color = 2'b11;
      12'h747: color = 2'b11;
      12'h748: color = 2'b11;
      12'h749: color = 2'b11;
      12'h74a: color = 2'b11;
      12'h74b: color = 2'b11;
      12'h74c: color = 2'b11;
      12'h74d: color = 2'b11;
      12'h74e: color = 2'b11;
      12'h74f: color = 2'b11;
      12'h750: color = 2'b01;
      12'h751: color = 2'b01;
      12'h752: color = 2'b00;
      12'h753: color = 2'b00;
      12'h754: color = 2'b00;
      12'h755: color = 2'b00;
      12'h756: color = 2'b00;
      12'h757: color = 2'b00;
      12'h758: color = 2'b00;
      12'h759: color = 2'b00;
      12'h75a: color = 2'b00;
      12'h75b: color = 2'b00;
      12'h75c: color = 2'b00;
      12'h75d: color = 2'b00;
      12'h75e: color = 2'b00;
      12'h75f: color = 2'b00;
      12'h760: color = 2'b00;
      12'h761: color = 2'b00;
      12'h762: color = 2'b01;
      12'h763: color = 2'b01;
      12'h764: color = 2'b01;
      12'h765: color = 2'b00;
      12'h766: color = 2'b00;
      12'h767: color = 2'b10;
      12'h768: color = 2'b10;
      12'h769: color = 2'b11;
      12'h76a: color = 2'b11;
      12'h76b: color = 2'b11;
      12'h76c: color = 2'b11;
      12'h76d: color = 2'b11;
      12'h76e: color = 2'b00;
      12'h76f: color = 2'b00;
      12'h770: color = 2'b11;
      12'h771: color = 2'b11;
      12'h772: color = 2'b11;
      12'h773: color = 2'b11;
      12'h774: color = 2'b11;
      12'h775: color = 2'b11;
      12'h776: color = 2'b11;
      12'h777: color = 2'b11;
      12'h778: color = 2'b11;
      12'h779: color = 2'b11;
      12'h77a: color = 2'b11;
      12'h77b: color = 2'b11;
      12'h77c: color = 2'b11;
      12'h77d: color = 2'b11;
      12'h77e: color = 2'b11;
      12'h77f: color = 2'b11;
      12'h780: color = 2'b11;
      12'h781: color = 2'b11;
      12'h782: color = 2'b11;
      12'h783: color = 2'b11;
      12'h784: color = 2'b11;
      12'h785: color = 2'b11;
      12'h786: color = 2'b11;
      12'h787: color = 2'b11;
      12'h788: color = 2'b11;
      12'h789: color = 2'b11;
      12'h78a: color = 2'b11;
      12'h78b: color = 2'b11;
      12'h78c: color = 2'b11;
      12'h78d: color = 2'b11;
      12'h78e: color = 2'b11;
      12'h78f: color = 2'b11;
      12'h790: color = 2'b01;
      12'h791: color = 2'b01;
      12'h792: color = 2'b00;
      12'h793: color = 2'b00;
      12'h794: color = 2'b00;
      12'h795: color = 2'b00;
      12'h796: color = 2'b00;
      12'h797: color = 2'b00;
      12'h798: color = 2'b00;
      12'h799: color = 2'b00;
      12'h79a: color = 2'b00;
      12'h79b: color = 2'b00;
      12'h79c: color = 2'b00;
      12'h79d: color = 2'b00;
      12'h79e: color = 2'b00;
      12'h79f: color = 2'b00;
      12'h7a0: color = 2'b00;
      12'h7a1: color = 2'b00;
      12'h7a2: color = 2'b01;
      12'h7a3: color = 2'b01;
      12'h7a4: color = 2'b01;
      12'h7a5: color = 2'b00;
      12'h7a6: color = 2'b00;
      12'h7a7: color = 2'b10;
      12'h7a8: color = 2'b10;
      12'h7a9: color = 2'b11;
      12'h7aa: color = 2'b11;
      12'h7ab: color = 2'b11;
      12'h7ac: color = 2'b11;
      12'h7ad: color = 2'b11;
      12'h7ae: color = 2'b00;
      12'h7af: color = 2'b00;
      12'h7b0: color = 2'b11;
      12'h7b1: color = 2'b11;
      12'h7b2: color = 2'b11;
      12'h7b3: color = 2'b11;
      12'h7b4: color = 2'b11;
      12'h7b5: color = 2'b11;
      12'h7b6: color = 2'b11;
      12'h7b7: color = 2'b11;
      12'h7b8: color = 2'b11;
      12'h7b9: color = 2'b11;
      12'h7ba: color = 2'b11;
      12'h7bb: color = 2'b11;
      12'h7bc: color = 2'b11;
      12'h7bd: color = 2'b11;
      12'h7be: color = 2'b11;
      12'h7bf: color = 2'b11;
      12'h7c0: color = 2'b11;
      12'h7c1: color = 2'b11;
      12'h7c2: color = 2'b11;
      12'h7c3: color = 2'b11;
      12'h7c4: color = 2'b11;
      12'h7c5: color = 2'b11;
      12'h7c6: color = 2'b11;
      12'h7c7: color = 2'b11;
      12'h7c8: color = 2'b11;
      12'h7c9: color = 2'b11;
      12'h7ca: color = 2'b11;
      12'h7cb: color = 2'b11;
      12'h7cc: color = 2'b11;
      12'h7cd: color = 2'b11;
      12'h7ce: color = 2'b11;
      12'h7cf: color = 2'b11;
      12'h7d0: color = 2'b01;
      12'h7d1: color = 2'b01;
      12'h7d2: color = 2'b00;
      12'h7d3: color = 2'b00;
      12'h7d4: color = 2'b00;
      12'h7d5: color = 2'b00;
      12'h7d6: color = 2'b00;
      12'h7d7: color = 2'b00;
      12'h7d8: color = 2'b00;
      12'h7d9: color = 2'b00;
      12'h7da: color = 2'b00;
      12'h7db: color = 2'b00;
      12'h7dc: color = 2'b00;
      12'h7dd: color = 2'b00;
      12'h7de: color = 2'b00;
      12'h7df: color = 2'b00;
      12'h7e0: color = 2'b00;
      12'h7e1: color = 2'b00;
      12'h7e2: color = 2'b01;
      12'h7e3: color = 2'b01;
      12'h7e4: color = 2'b01;
      12'h7e5: color = 2'b00;
      12'h7e6: color = 2'b00;
      12'h7e7: color = 2'b10;
      12'h7e8: color = 2'b10;
      12'h7e9: color = 2'b11;
      12'h7ea: color = 2'b11;
      12'h7eb: color = 2'b11;
      12'h7ec: color = 2'b11;
      12'h7ed: color = 2'b11;
      12'h7ee: color = 2'b00;
      12'h7ef: color = 2'b00;
      12'h7f0: color = 2'b11;
      12'h7f1: color = 2'b11;
      12'h7f2: color = 2'b11;
      12'h7f3: color = 2'b11;
      12'h7f4: color = 2'b11;
      12'h7f5: color = 2'b11;
      12'h7f6: color = 2'b11;
      12'h7f7: color = 2'b11;
      12'h7f8: color = 2'b11;
      12'h7f9: color = 2'b11;
      12'h7fa: color = 2'b11;
      12'h7fb: color = 2'b11;
      12'h7fc: color = 2'b11;
      12'h7fd: color = 2'b11;
      12'h7fe: color = 2'b11;
      12'h7ff: color = 2'b11;
      12'h800: color = 2'b11;
      12'h801: color = 2'b11;
      12'h802: color = 2'b11;
      12'h803: color = 2'b11;
      12'h804: color = 2'b11;
      12'h805: color = 2'b11;
      12'h806: color = 2'b11;
      12'h807: color = 2'b11;
      12'h808: color = 2'b11;
      12'h809: color = 2'b11;
      12'h80a: color = 2'b11;
      12'h80b: color = 2'b11;
      12'h80c: color = 2'b11;
      12'h80d: color = 2'b11;
      12'h80e: color = 2'b11;
      12'h80f: color = 2'b11;
      12'h810: color = 2'b11;
      12'h811: color = 2'b11;
      12'h812: color = 2'b01;
      12'h813: color = 2'b01;
      12'h814: color = 2'b01;
      12'h815: color = 2'b00;
      12'h816: color = 2'b00;
      12'h817: color = 2'b00;
      12'h818: color = 2'b00;
      12'h819: color = 2'b00;
      12'h81a: color = 2'b00;
      12'h81b: color = 2'b00;
      12'h81c: color = 2'b00;
      12'h81d: color = 2'b00;
      12'h81e: color = 2'b01;
      12'h81f: color = 2'b01;
      12'h820: color = 2'b10;
      12'h821: color = 2'b10;
      12'h822: color = 2'b10;
      12'h823: color = 2'b10;
      12'h824: color = 2'b10;
      12'h825: color = 2'b10;
      12'h826: color = 2'b10;
      12'h827: color = 2'b10;
      12'h828: color = 2'b10;
      12'h829: color = 2'b10;
      12'h82a: color = 2'b10;
      12'h82b: color = 2'b00;
      12'h82c: color = 2'b00;
      12'h82d: color = 2'b00;
      12'h82e: color = 2'b11;
      12'h82f: color = 2'b11;
      12'h830: color = 2'b11;
      12'h831: color = 2'b11;
      12'h832: color = 2'b11;
      12'h833: color = 2'b11;
      12'h834: color = 2'b11;
      12'h835: color = 2'b11;
      12'h836: color = 2'b11;
      12'h837: color = 2'b11;
      12'h838: color = 2'b11;
      12'h839: color = 2'b11;
      12'h83a: color = 2'b11;
      12'h83b: color = 2'b11;
      12'h83c: color = 2'b11;
      12'h83d: color = 2'b11;
      12'h83e: color = 2'b11;
      12'h83f: color = 2'b11;
      12'h840: color = 2'b11;
      12'h841: color = 2'b11;
      12'h842: color = 2'b11;
      12'h843: color = 2'b11;
      12'h844: color = 2'b11;
      12'h845: color = 2'b11;
      12'h846: color = 2'b11;
      12'h847: color = 2'b11;
      12'h848: color = 2'b11;
      12'h849: color = 2'b11;
      12'h84a: color = 2'b11;
      12'h84b: color = 2'b11;
      12'h84c: color = 2'b11;
      12'h84d: color = 2'b11;
      12'h84e: color = 2'b11;
      12'h84f: color = 2'b11;
      12'h850: color = 2'b11;
      12'h851: color = 2'b11;
      12'h852: color = 2'b01;
      12'h853: color = 2'b01;
      12'h854: color = 2'b01;
      12'h855: color = 2'b00;
      12'h856: color = 2'b00;
      12'h857: color = 2'b00;
      12'h858: color = 2'b00;
      12'h859: color = 2'b00;
      12'h85a: color = 2'b00;
      12'h85b: color = 2'b00;
      12'h85c: color = 2'b00;
      12'h85d: color = 2'b00;
      12'h85e: color = 2'b01;
      12'h85f: color = 2'b01;
      12'h860: color = 2'b10;
      12'h861: color = 2'b10;
      12'h862: color = 2'b10;
      12'h863: color = 2'b10;
      12'h864: color = 2'b10;
      12'h865: color = 2'b10;
      12'h866: color = 2'b10;
      12'h867: color = 2'b10;
      12'h868: color = 2'b10;
      12'h869: color = 2'b10;
      12'h86a: color = 2'b10;
      12'h86b: color = 2'b00;
      12'h86c: color = 2'b00;
      12'h86d: color = 2'b00;
      12'h86e: color = 2'b11;
      12'h86f: color = 2'b11;
      12'h870: color = 2'b11;
      12'h871: color = 2'b11;
      12'h872: color = 2'b11;
      12'h873: color = 2'b11;
      12'h874: color = 2'b11;
      12'h875: color = 2'b11;
      12'h876: color = 2'b11;
      12'h877: color = 2'b11;
      12'h878: color = 2'b11;
      12'h879: color = 2'b11;
      12'h87a: color = 2'b11;
      12'h87b: color = 2'b11;
      12'h87c: color = 2'b11;
      12'h87d: color = 2'b11;
      12'h87e: color = 2'b11;
      12'h87f: color = 2'b11;
      12'h880: color = 2'b11;
      12'h881: color = 2'b11;
      12'h882: color = 2'b11;
      12'h883: color = 2'b11;
      12'h884: color = 2'b11;
      12'h885: color = 2'b11;
      12'h886: color = 2'b11;
      12'h887: color = 2'b11;
      12'h888: color = 2'b11;
      12'h889: color = 2'b11;
      12'h88a: color = 2'b11;
      12'h88b: color = 2'b01;
      12'h88c: color = 2'b01;
      12'h88d: color = 2'b01;
      12'h88e: color = 2'b00;
      12'h88f: color = 2'b00;
      12'h890: color = 2'b00;
      12'h891: color = 2'b00;
      12'h892: color = 2'b00;
      12'h893: color = 2'b00;
      12'h894: color = 2'b00;
      12'h895: color = 2'b00;
      12'h896: color = 2'b00;
      12'h897: color = 2'b01;
      12'h898: color = 2'b01;
      12'h899: color = 2'b01;
      12'h89a: color = 2'b01;
      12'h89b: color = 2'b01;
      12'h89c: color = 2'b01;
      12'h89d: color = 2'b01;
      12'h89e: color = 2'b00;
      12'h89f: color = 2'b00;
      12'h8a0: color = 2'b00;
      12'h8a1: color = 2'b00;
      12'h8a2: color = 2'b01;
      12'h8a3: color = 2'b01;
      12'h8a4: color = 2'b01;
      12'h8a5: color = 2'b01;
      12'h8a6: color = 2'b01;
      12'h8a7: color = 2'b00;
      12'h8a8: color = 2'b00;
      12'h8a9: color = 2'b01;
      12'h8aa: color = 2'b01;
      12'h8ab: color = 2'b11;
      12'h8ac: color = 2'b11;
      12'h8ad: color = 2'b11;
      12'h8ae: color = 2'b11;
      12'h8af: color = 2'b11;
      12'h8b0: color = 2'b11;
      12'h8b1: color = 2'b11;
      12'h8b2: color = 2'b11;
      12'h8b3: color = 2'b11;
      12'h8b4: color = 2'b11;
      12'h8b5: color = 2'b11;
      12'h8b6: color = 2'b11;
      12'h8b7: color = 2'b11;
      12'h8b8: color = 2'b11;
      12'h8b9: color = 2'b11;
      12'h8ba: color = 2'b11;
      12'h8bb: color = 2'b11;
      12'h8bc: color = 2'b11;
      12'h8bd: color = 2'b11;
      12'h8be: color = 2'b11;
      12'h8bf: color = 2'b11;
      12'h8c0: color = 2'b11;
      12'h8c1: color = 2'b11;
      12'h8c2: color = 2'b11;
      12'h8c3: color = 2'b11;
      12'h8c4: color = 2'b11;
      12'h8c5: color = 2'b11;
      12'h8c6: color = 2'b11;
      12'h8c7: color = 2'b11;
      12'h8c8: color = 2'b11;
      12'h8c9: color = 2'b11;
      12'h8ca: color = 2'b11;
      12'h8cb: color = 2'b01;
      12'h8cc: color = 2'b01;
      12'h8cd: color = 2'b01;
      12'h8ce: color = 2'b00;
      12'h8cf: color = 2'b00;
      12'h8d0: color = 2'b00;
      12'h8d1: color = 2'b00;
      12'h8d2: color = 2'b00;
      12'h8d3: color = 2'b00;
      12'h8d4: color = 2'b00;
      12'h8d5: color = 2'b00;
      12'h8d6: color = 2'b00;
      12'h8d7: color = 2'b01;
      12'h8d8: color = 2'b01;
      12'h8d9: color = 2'b01;
      12'h8da: color = 2'b01;
      12'h8db: color = 2'b01;
      12'h8dc: color = 2'b01;
      12'h8dd: color = 2'b01;
      12'h8de: color = 2'b00;
      12'h8df: color = 2'b00;
      12'h8e0: color = 2'b00;
      12'h8e1: color = 2'b00;
      12'h8e2: color = 2'b01;
      12'h8e3: color = 2'b01;
      12'h8e4: color = 2'b01;
      12'h8e5: color = 2'b01;
      12'h8e6: color = 2'b01;
      12'h8e7: color = 2'b00;
      12'h8e8: color = 2'b00;
      12'h8e9: color = 2'b01;
      12'h8ea: color = 2'b01;
      12'h8eb: color = 2'b11;
      12'h8ec: color = 2'b11;
      12'h8ed: color = 2'b11;
      12'h8ee: color = 2'b11;
      12'h8ef: color = 2'b11;
      12'h8f0: color = 2'b11;
      12'h8f1: color = 2'b11;
      12'h8f2: color = 2'b11;
      12'h8f3: color = 2'b11;
      12'h8f4: color = 2'b11;
      12'h8f5: color = 2'b11;
      12'h8f6: color = 2'b11;
      12'h8f7: color = 2'b11;
      12'h8f8: color = 2'b11;
      12'h8f9: color = 2'b11;
      12'h8fa: color = 2'b11;
      12'h8fb: color = 2'b11;
      12'h8fc: color = 2'b11;
      12'h8fd: color = 2'b11;
      12'h8fe: color = 2'b11;
      12'h8ff: color = 2'b11;
      12'h900: color = 2'b11;
      12'h901: color = 2'b11;
      12'h902: color = 2'b11;
      12'h903: color = 2'b11;
      12'h904: color = 2'b11;
      12'h905: color = 2'b11;
      12'h906: color = 2'b11;
      12'h907: color = 2'b01;
      12'h908: color = 2'b01;
      12'h909: color = 2'b00;
      12'h90a: color = 2'b00;
      12'h90b: color = 2'b10;
      12'h90c: color = 2'b10;
      12'h90d: color = 2'b10;
      12'h90e: color = 2'b10;
      12'h90f: color = 2'b10;
      12'h910: color = 2'b10;
      12'h911: color = 2'b10;
      12'h912: color = 2'b10;
      12'h913: color = 2'b10;
      12'h914: color = 2'b10;
      12'h915: color = 2'b10;
      12'h916: color = 2'b10;
      12'h917: color = 2'b00;
      12'h918: color = 2'b00;
      12'h919: color = 2'b00;
      12'h91a: color = 2'b00;
      12'h91b: color = 2'b00;
      12'h91c: color = 2'b00;
      12'h91d: color = 2'b00;
      12'h91e: color = 2'b01;
      12'h91f: color = 2'b01;
      12'h920: color = 2'b01;
      12'h921: color = 2'b01;
      12'h922: color = 2'b00;
      12'h923: color = 2'b00;
      12'h924: color = 2'b00;
      12'h925: color = 2'b00;
      12'h926: color = 2'b00;
      12'h927: color = 2'b11;
      12'h928: color = 2'b11;
      12'h929: color = 2'b11;
      12'h92a: color = 2'b11;
      12'h92b: color = 2'b11;
      12'h92c: color = 2'b11;
      12'h92d: color = 2'b11;
      12'h92e: color = 2'b11;
      12'h92f: color = 2'b11;
      12'h930: color = 2'b11;
      12'h931: color = 2'b11;
      12'h932: color = 2'b11;
      12'h933: color = 2'b11;
      12'h934: color = 2'b11;
      12'h935: color = 2'b11;
      12'h936: color = 2'b11;
      12'h937: color = 2'b11;
      12'h938: color = 2'b11;
      12'h939: color = 2'b11;
      12'h93a: color = 2'b11;
      12'h93b: color = 2'b11;
      12'h93c: color = 2'b11;
      12'h93d: color = 2'b11;
      12'h93e: color = 2'b11;
      12'h93f: color = 2'b11;
      12'h940: color = 2'b11;
      12'h941: color = 2'b11;
      12'h942: color = 2'b11;
      12'h943: color = 2'b11;
      12'h944: color = 2'b11;
      12'h945: color = 2'b11;
      12'h946: color = 2'b11;
      12'h947: color = 2'b01;
      12'h948: color = 2'b01;
      12'h949: color = 2'b00;
      12'h94a: color = 2'b00;
      12'h94b: color = 2'b10;
      12'h94c: color = 2'b10;
      12'h94d: color = 2'b10;
      12'h94e: color = 2'b10;
      12'h94f: color = 2'b10;
      12'h950: color = 2'b10;
      12'h951: color = 2'b10;
      12'h952: color = 2'b10;
      12'h953: color = 2'b10;
      12'h954: color = 2'b10;
      12'h955: color = 2'b10;
      12'h956: color = 2'b10;
      12'h957: color = 2'b00;
      12'h958: color = 2'b00;
      12'h959: color = 2'b00;
      12'h95a: color = 2'b00;
      12'h95b: color = 2'b00;
      12'h95c: color = 2'b00;
      12'h95d: color = 2'b00;
      12'h95e: color = 2'b01;
      12'h95f: color = 2'b01;
      12'h960: color = 2'b01;
      12'h961: color = 2'b01;
      12'h962: color = 2'b00;
      12'h963: color = 2'b00;
      12'h964: color = 2'b00;
      12'h965: color = 2'b00;
      12'h966: color = 2'b00;
      12'h967: color = 2'b11;
      12'h968: color = 2'b11;
      12'h969: color = 2'b11;
      12'h96a: color = 2'b11;
      12'h96b: color = 2'b11;
      12'h96c: color = 2'b11;
      12'h96d: color = 2'b11;
      12'h96e: color = 2'b11;
      12'h96f: color = 2'b11;
      12'h970: color = 2'b11;
      12'h971: color = 2'b11;
      12'h972: color = 2'b11;
      12'h973: color = 2'b11;
      12'h974: color = 2'b11;
      12'h975: color = 2'b11;
      12'h976: color = 2'b11;
      12'h977: color = 2'b11;
      12'h978: color = 2'b11;
      12'h979: color = 2'b11;
      12'h97a: color = 2'b11;
      12'h97b: color = 2'b11;
      12'h97c: color = 2'b11;
      12'h97d: color = 2'b11;
      12'h97e: color = 2'b11;
      12'h97f: color = 2'b11;
      12'h980: color = 2'b11;
      12'h981: color = 2'b11;
      12'h982: color = 2'b11;
      12'h983: color = 2'b11;
      12'h984: color = 2'b11;
      12'h985: color = 2'b11;
      12'h986: color = 2'b11;
      12'h987: color = 2'b01;
      12'h988: color = 2'b01;
      12'h989: color = 2'b00;
      12'h98a: color = 2'b00;
      12'h98b: color = 2'b10;
      12'h98c: color = 2'b10;
      12'h98d: color = 2'b10;
      12'h98e: color = 2'b10;
      12'h98f: color = 2'b10;
      12'h990: color = 2'b10;
      12'h991: color = 2'b10;
      12'h992: color = 2'b10;
      12'h993: color = 2'b10;
      12'h994: color = 2'b10;
      12'h995: color = 2'b10;
      12'h996: color = 2'b10;
      12'h997: color = 2'b00;
      12'h998: color = 2'b00;
      12'h999: color = 2'b00;
      12'h99a: color = 2'b00;
      12'h99b: color = 2'b00;
      12'h99c: color = 2'b00;
      12'h99d: color = 2'b00;
      12'h99e: color = 2'b01;
      12'h99f: color = 2'b01;
      12'h9a0: color = 2'b01;
      12'h9a1: color = 2'b01;
      12'h9a2: color = 2'b00;
      12'h9a3: color = 2'b00;
      12'h9a4: color = 2'b00;
      12'h9a5: color = 2'b00;
      12'h9a6: color = 2'b00;
      12'h9a7: color = 2'b11;
      12'h9a8: color = 2'b11;
      12'h9a9: color = 2'b11;
      12'h9aa: color = 2'b11;
      12'h9ab: color = 2'b11;
      12'h9ac: color = 2'b11;
      12'h9ad: color = 2'b11;
      12'h9ae: color = 2'b11;
      12'h9af: color = 2'b11;
      12'h9b0: color = 2'b11;
      12'h9b1: color = 2'b11;
      12'h9b2: color = 2'b11;
      12'h9b3: color = 2'b11;
      12'h9b4: color = 2'b11;
      12'h9b5: color = 2'b11;
      12'h9b6: color = 2'b11;
      12'h9b7: color = 2'b11;
      12'h9b8: color = 2'b11;
      12'h9b9: color = 2'b11;
      12'h9ba: color = 2'b11;
      12'h9bb: color = 2'b11;
      12'h9bc: color = 2'b11;
      12'h9bd: color = 2'b11;
      12'h9be: color = 2'b11;
      12'h9bf: color = 2'b11;
      12'h9c0: color = 2'b11;
      12'h9c1: color = 2'b11;
      12'h9c2: color = 2'b11;
      12'h9c3: color = 2'b11;
      12'h9c4: color = 2'b11;
      12'h9c5: color = 2'b01;
      12'h9c6: color = 2'b01;
      12'h9c7: color = 2'b10;
      12'h9c8: color = 2'b10;
      12'h9c9: color = 2'b01;
      12'h9ca: color = 2'b01;
      12'h9cb: color = 2'b10;
      12'h9cc: color = 2'b10;
      12'h9cd: color = 2'b10;
      12'h9ce: color = 2'b10;
      12'h9cf: color = 2'b10;
      12'h9d0: color = 2'b10;
      12'h9d1: color = 2'b10;
      12'h9d2: color = 2'b10;
      12'h9d3: color = 2'b10;
      12'h9d4: color = 2'b10;
      12'h9d5: color = 2'b10;
      12'h9d6: color = 2'b10;
      12'h9d7: color = 2'b10;
      12'h9d8: color = 2'b10;
      12'h9d9: color = 2'b10;
      12'h9da: color = 2'b10;
      12'h9db: color = 2'b00;
      12'h9dc: color = 2'b00;
      12'h9dd: color = 2'b00;
      12'h9de: color = 2'b00;
      12'h9df: color = 2'b00;
      12'h9e0: color = 2'b01;
      12'h9e1: color = 2'b01;
      12'h9e2: color = 2'b00;
      12'h9e3: color = 2'b00;
      12'h9e4: color = 2'b00;
      12'h9e5: color = 2'b11;
      12'h9e6: color = 2'b11;
      12'h9e7: color = 2'b00;
      12'h9e8: color = 2'b00;
      12'h9e9: color = 2'b01;
      12'h9ea: color = 2'b01;
      12'h9eb: color = 2'b11;
      12'h9ec: color = 2'b11;
      12'h9ed: color = 2'b11;
      12'h9ee: color = 2'b11;
      12'h9ef: color = 2'b11;
      12'h9f0: color = 2'b11;
      12'h9f1: color = 2'b11;
      12'h9f2: color = 2'b11;
      12'h9f3: color = 2'b11;
      12'h9f4: color = 2'b11;
      12'h9f5: color = 2'b11;
      12'h9f6: color = 2'b11;
      12'h9f7: color = 2'b11;
      12'h9f8: color = 2'b11;
      12'h9f9: color = 2'b11;
      12'h9fa: color = 2'b11;
      12'h9fb: color = 2'b11;
      12'h9fc: color = 2'b11;
      12'h9fd: color = 2'b11;
      12'h9fe: color = 2'b11;
      12'h9ff: color = 2'b11;
      12'ha00: color = 2'b11;
      12'ha01: color = 2'b11;
      12'ha02: color = 2'b11;
      12'ha03: color = 2'b11;
      12'ha04: color = 2'b11;
      12'ha05: color = 2'b01;
      12'ha06: color = 2'b01;
      12'ha07: color = 2'b10;
      12'ha08: color = 2'b10;
      12'ha09: color = 2'b01;
      12'ha0a: color = 2'b01;
      12'ha0b: color = 2'b10;
      12'ha0c: color = 2'b10;
      12'ha0d: color = 2'b10;
      12'ha0e: color = 2'b10;
      12'ha0f: color = 2'b10;
      12'ha10: color = 2'b10;
      12'ha11: color = 2'b10;
      12'ha12: color = 2'b10;
      12'ha13: color = 2'b10;
      12'ha14: color = 2'b10;
      12'ha15: color = 2'b10;
      12'ha16: color = 2'b10;
      12'ha17: color = 2'b10;
      12'ha18: color = 2'b10;
      12'ha19: color = 2'b10;
      12'ha1a: color = 2'b10;
      12'ha1b: color = 2'b00;
      12'ha1c: color = 2'b00;
      12'ha1d: color = 2'b00;
      12'ha1e: color = 2'b00;
      12'ha1f: color = 2'b00;
      12'ha20: color = 2'b01;
      12'ha21: color = 2'b01;
      12'ha22: color = 2'b00;
      12'ha23: color = 2'b00;
      12'ha24: color = 2'b00;
      12'ha25: color = 2'b11;
      12'ha26: color = 2'b11;
      12'ha27: color = 2'b00;
      12'ha28: color = 2'b00;
      12'ha29: color = 2'b01;
      12'ha2a: color = 2'b01;
      12'ha2b: color = 2'b11;
      12'ha2c: color = 2'b11;
      12'ha2d: color = 2'b11;
      12'ha2e: color = 2'b11;
      12'ha2f: color = 2'b11;
      12'ha30: color = 2'b11;
      12'ha31: color = 2'b11;
      12'ha32: color = 2'b11;
      12'ha33: color = 2'b11;
      12'ha34: color = 2'b11;
      12'ha35: color = 2'b11;
      12'ha36: color = 2'b11;
      12'ha37: color = 2'b11;
      12'ha38: color = 2'b11;
      12'ha39: color = 2'b11;
      12'ha3a: color = 2'b11;
      12'ha3b: color = 2'b11;
      12'ha3c: color = 2'b11;
      12'ha3d: color = 2'b11;
      12'ha3e: color = 2'b11;
      12'ha3f: color = 2'b11;
      12'ha40: color = 2'b11;
      12'ha41: color = 2'b11;
      12'ha42: color = 2'b11;
      12'ha43: color = 2'b11;
      12'ha44: color = 2'b11;
      12'ha45: color = 2'b00;
      12'ha46: color = 2'b00;
      12'ha47: color = 2'b01;
      12'ha48: color = 2'b01;
      12'ha49: color = 2'b10;
      12'ha4a: color = 2'b10;
      12'ha4b: color = 2'b01;
      12'ha4c: color = 2'b01;
      12'ha4d: color = 2'b01;
      12'ha4e: color = 2'b10;
      12'ha4f: color = 2'b10;
      12'ha50: color = 2'b01;
      12'ha51: color = 2'b01;
      12'ha52: color = 2'b10;
      12'ha53: color = 2'b10;
      12'ha54: color = 2'b10;
      12'ha55: color = 2'b01;
      12'ha56: color = 2'b01;
      12'ha57: color = 2'b10;
      12'ha58: color = 2'b10;
      12'ha59: color = 2'b00;
      12'ha5a: color = 2'b00;
      12'ha5b: color = 2'b00;
      12'ha5c: color = 2'b00;
      12'ha5d: color = 2'b00;
      12'ha5e: color = 2'b01;
      12'ha5f: color = 2'b01;
      12'ha60: color = 2'b00;
      12'ha61: color = 2'b00;
      12'ha62: color = 2'b10;
      12'ha63: color = 2'b10;
      12'ha64: color = 2'b10;
      12'ha65: color = 2'b11;
      12'ha66: color = 2'b11;
      12'ha67: color = 2'b11;
      12'ha68: color = 2'b11;
      12'ha69: color = 2'b11;
      12'ha6a: color = 2'b11;
      12'ha6b: color = 2'b00;
      12'ha6c: color = 2'b00;
      12'ha6d: color = 2'b00;
      12'ha6e: color = 2'b11;
      12'ha6f: color = 2'b11;
      12'ha70: color = 2'b11;
      12'ha71: color = 2'b11;
      12'ha72: color = 2'b11;
      12'ha73: color = 2'b11;
      12'ha74: color = 2'b11;
      12'ha75: color = 2'b11;
      12'ha76: color = 2'b11;
      12'ha77: color = 2'b11;
      12'ha78: color = 2'b11;
      12'ha79: color = 2'b11;
      12'ha7a: color = 2'b11;
      12'ha7b: color = 2'b11;
      12'ha7c: color = 2'b11;
      12'ha7d: color = 2'b11;
      12'ha7e: color = 2'b11;
      12'ha7f: color = 2'b11;
      12'ha80: color = 2'b11;
      12'ha81: color = 2'b11;
      12'ha82: color = 2'b11;
      12'ha83: color = 2'b11;
      12'ha84: color = 2'b11;
      12'ha85: color = 2'b00;
      12'ha86: color = 2'b00;
      12'ha87: color = 2'b01;
      12'ha88: color = 2'b01;
      12'ha89: color = 2'b10;
      12'ha8a: color = 2'b10;
      12'ha8b: color = 2'b01;
      12'ha8c: color = 2'b01;
      12'ha8d: color = 2'b01;
      12'ha8e: color = 2'b10;
      12'ha8f: color = 2'b10;
      12'ha90: color = 2'b01;
      12'ha91: color = 2'b01;
      12'ha92: color = 2'b10;
      12'ha93: color = 2'b10;
      12'ha94: color = 2'b10;
      12'ha95: color = 2'b01;
      12'ha96: color = 2'b01;
      12'ha97: color = 2'b10;
      12'ha98: color = 2'b10;
      12'ha99: color = 2'b00;
      12'ha9a: color = 2'b00;
      12'ha9b: color = 2'b00;
      12'ha9c: color = 2'b00;
      12'ha9d: color = 2'b00;
      12'ha9e: color = 2'b01;
      12'ha9f: color = 2'b01;
      12'haa0: color = 2'b00;
      12'haa1: color = 2'b00;
      12'haa2: color = 2'b10;
      12'haa3: color = 2'b10;
      12'haa4: color = 2'b10;
      12'haa5: color = 2'b11;
      12'haa6: color = 2'b11;
      12'haa7: color = 2'b11;
      12'haa8: color = 2'b11;
      12'haa9: color = 2'b11;
      12'haaa: color = 2'b11;
      12'haab: color = 2'b00;
      12'haac: color = 2'b00;
      12'haad: color = 2'b00;
      12'haae: color = 2'b11;
      12'haaf: color = 2'b11;
      12'hab0: color = 2'b11;
      12'hab1: color = 2'b11;
      12'hab2: color = 2'b11;
      12'hab3: color = 2'b11;
      12'hab4: color = 2'b11;
      12'hab5: color = 2'b11;
      12'hab6: color = 2'b11;
      12'hab7: color = 2'b11;
      12'hab8: color = 2'b11;
      12'hab9: color = 2'b11;
      12'haba: color = 2'b11;
      12'habb: color = 2'b11;
      12'habc: color = 2'b11;
      12'habd: color = 2'b11;
      12'habe: color = 2'b11;
      12'habf: color = 2'b11;
      12'hac0: color = 2'b11;
      12'hac1: color = 2'b11;
      12'hac2: color = 2'b00;
      12'hac3: color = 2'b00;
      12'hac4: color = 2'b00;
      12'hac5: color = 2'b01;
      12'hac6: color = 2'b01;
      12'hac7: color = 2'b01;
      12'hac8: color = 2'b01;
      12'hac9: color = 2'b00;
      12'haca: color = 2'b00;
      12'hacb: color = 2'b00;
      12'hacc: color = 2'b00;
      12'hacd: color = 2'b00;
      12'hace: color = 2'b01;
      12'hacf: color = 2'b01;
      12'had0: color = 2'b10;
      12'had1: color = 2'b10;
      12'had2: color = 2'b01;
      12'had3: color = 2'b01;
      12'had4: color = 2'b01;
      12'had5: color = 2'b10;
      12'had6: color = 2'b10;
      12'had7: color = 2'b00;
      12'had8: color = 2'b00;
      12'had9: color = 2'b01;
      12'hada: color = 2'b01;
      12'hadb: color = 2'b01;
      12'hadc: color = 2'b01;
      12'hadd: color = 2'b01;
      12'hade: color = 2'b01;
      12'hadf: color = 2'b01;
      12'hae0: color = 2'b00;
      12'hae1: color = 2'b00;
      12'hae2: color = 2'b10;
      12'hae3: color = 2'b10;
      12'hae4: color = 2'b10;
      12'hae5: color = 2'b11;
      12'hae6: color = 2'b11;
      12'hae7: color = 2'b11;
      12'hae8: color = 2'b11;
      12'hae9: color = 2'b00;
      12'haea: color = 2'b00;
      12'haeb: color = 2'b11;
      12'haec: color = 2'b11;
      12'haed: color = 2'b11;
      12'haee: color = 2'b00;
      12'haef: color = 2'b00;
      12'haf0: color = 2'b11;
      12'haf1: color = 2'b11;
      12'haf2: color = 2'b11;
      12'haf3: color = 2'b11;
      12'haf4: color = 2'b11;
      12'haf5: color = 2'b00;
      12'haf6: color = 2'b00;
      12'haf7: color = 2'b00;
      12'haf8: color = 2'b00;
      12'haf9: color = 2'b01;
      12'hafa: color = 2'b01;
      12'hafb: color = 2'b11;
      12'hafc: color = 2'b11;
      12'hafd: color = 2'b11;
      12'hafe: color = 2'b11;
      12'haff: color = 2'b11;
      12'hb00: color = 2'b11;
      12'hb01: color = 2'b11;
      12'hb02: color = 2'b00;
      12'hb03: color = 2'b00;
      12'hb04: color = 2'b00;
      12'hb05: color = 2'b01;
      12'hb06: color = 2'b01;
      12'hb07: color = 2'b01;
      12'hb08: color = 2'b01;
      12'hb09: color = 2'b00;
      12'hb0a: color = 2'b00;
      12'hb0b: color = 2'b00;
      12'hb0c: color = 2'b00;
      12'hb0d: color = 2'b00;
      12'hb0e: color = 2'b01;
      12'hb0f: color = 2'b01;
      12'hb10: color = 2'b10;
      12'hb11: color = 2'b10;
      12'hb12: color = 2'b01;
      12'hb13: color = 2'b01;
      12'hb14: color = 2'b01;
      12'hb15: color = 2'b10;
      12'hb16: color = 2'b10;
      12'hb17: color = 2'b00;
      12'hb18: color = 2'b00;
      12'hb19: color = 2'b01;
      12'hb1a: color = 2'b01;
      12'hb1b: color = 2'b01;
      12'hb1c: color = 2'b01;
      12'hb1d: color = 2'b01;
      12'hb1e: color = 2'b01;
      12'hb1f: color = 2'b01;
      12'hb20: color = 2'b00;
      12'hb21: color = 2'b00;
      12'hb22: color = 2'b10;
      12'hb23: color = 2'b10;
      12'hb24: color = 2'b10;
      12'hb25: color = 2'b11;
      12'hb26: color = 2'b11;
      12'hb27: color = 2'b11;
      12'hb28: color = 2'b11;
      12'hb29: color = 2'b00;
      12'hb2a: color = 2'b00;
      12'hb2b: color = 2'b11;
      12'hb2c: color = 2'b11;
      12'hb2d: color = 2'b11;
      12'hb2e: color = 2'b00;
      12'hb2f: color = 2'b00;
      12'hb30: color = 2'b11;
      12'hb31: color = 2'b11;
      12'hb32: color = 2'b11;
      12'hb33: color = 2'b11;
      12'hb34: color = 2'b11;
      12'hb35: color = 2'b00;
      12'hb36: color = 2'b00;
      12'hb37: color = 2'b00;
      12'hb38: color = 2'b00;
      12'hb39: color = 2'b01;
      12'hb3a: color = 2'b01;
      12'hb3b: color = 2'b11;
      12'hb3c: color = 2'b11;
      12'hb3d: color = 2'b11;
      12'hb3e: color = 2'b11;
      12'hb3f: color = 2'b11;
      12'hb40: color = 2'b11;
      12'hb41: color = 2'b11;
      12'hb42: color = 2'b00;
      12'hb43: color = 2'b00;
      12'hb44: color = 2'b00;
      12'hb45: color = 2'b01;
      12'hb46: color = 2'b01;
      12'hb47: color = 2'b01;
      12'hb48: color = 2'b01;
      12'hb49: color = 2'b00;
      12'hb4a: color = 2'b00;
      12'hb4b: color = 2'b00;
      12'hb4c: color = 2'b00;
      12'hb4d: color = 2'b00;
      12'hb4e: color = 2'b01;
      12'hb4f: color = 2'b01;
      12'hb50: color = 2'b10;
      12'hb51: color = 2'b10;
      12'hb52: color = 2'b01;
      12'hb53: color = 2'b01;
      12'hb54: color = 2'b01;
      12'hb55: color = 2'b10;
      12'hb56: color = 2'b10;
      12'hb57: color = 2'b00;
      12'hb58: color = 2'b00;
      12'hb59: color = 2'b01;
      12'hb5a: color = 2'b01;
      12'hb5b: color = 2'b01;
      12'hb5c: color = 2'b01;
      12'hb5d: color = 2'b01;
      12'hb5e: color = 2'b01;
      12'hb5f: color = 2'b01;
      12'hb60: color = 2'b00;
      12'hb61: color = 2'b00;
      12'hb62: color = 2'b10;
      12'hb63: color = 2'b10;
      12'hb64: color = 2'b10;
      12'hb65: color = 2'b11;
      12'hb66: color = 2'b11;
      12'hb67: color = 2'b11;
      12'hb68: color = 2'b11;
      12'hb69: color = 2'b00;
      12'hb6a: color = 2'b00;
      12'hb6b: color = 2'b11;
      12'hb6c: color = 2'b11;
      12'hb6d: color = 2'b11;
      12'hb6e: color = 2'b00;
      12'hb6f: color = 2'b00;
      12'hb70: color = 2'b11;
      12'hb71: color = 2'b11;
      12'hb72: color = 2'b11;
      12'hb73: color = 2'b11;
      12'hb74: color = 2'b11;
      12'hb75: color = 2'b00;
      12'hb76: color = 2'b00;
      12'hb77: color = 2'b00;
      12'hb78: color = 2'b00;
      12'hb79: color = 2'b01;
      12'hb7a: color = 2'b01;
      12'hb7b: color = 2'b11;
      12'hb7c: color = 2'b11;
      12'hb7d: color = 2'b11;
      12'hb7e: color = 2'b11;
      12'hb7f: color = 2'b11;
      12'hb80: color = 2'b11;
      12'hb81: color = 2'b11;
      12'hb82: color = 2'b00;
      12'hb83: color = 2'b00;
      12'hb84: color = 2'b00;
      12'hb85: color = 2'b00;
      12'hb86: color = 2'b00;
      12'hb87: color = 2'b00;
      12'hb88: color = 2'b00;
      12'hb89: color = 2'b11;
      12'hb8a: color = 2'b11;
      12'hb8b: color = 2'b11;
      12'hb8c: color = 2'b11;
      12'hb8d: color = 2'b11;
      12'hb8e: color = 2'b00;
      12'hb8f: color = 2'b00;
      12'hb90: color = 2'b01;
      12'hb91: color = 2'b01;
      12'hb92: color = 2'b01;
      12'hb93: color = 2'b01;
      12'hb94: color = 2'b01;
      12'hb95: color = 2'b01;
      12'hb96: color = 2'b01;
      12'hb97: color = 2'b00;
      12'hb98: color = 2'b00;
      12'hb99: color = 2'b01;
      12'hb9a: color = 2'b01;
      12'hb9b: color = 2'b01;
      12'hb9c: color = 2'b01;
      12'hb9d: color = 2'b01;
      12'hb9e: color = 2'b01;
      12'hb9f: color = 2'b01;
      12'hba0: color = 2'b00;
      12'hba1: color = 2'b00;
      12'hba2: color = 2'b10;
      12'hba3: color = 2'b10;
      12'hba4: color = 2'b10;
      12'hba5: color = 2'b10;
      12'hba6: color = 2'b10;
      12'hba7: color = 2'b00;
      12'hba8: color = 2'b00;
      12'hba9: color = 2'b11;
      12'hbaa: color = 2'b11;
      12'hbab: color = 2'b11;
      12'hbac: color = 2'b11;
      12'hbad: color = 2'b11;
      12'hbae: color = 2'b11;
      12'hbaf: color = 2'b11;
      12'hbb0: color = 2'b00;
      12'hbb1: color = 2'b00;
      12'hbb2: color = 2'b00;
      12'hbb3: color = 2'b00;
      12'hbb4: color = 2'b00;
      12'hbb5: color = 2'b11;
      12'hbb6: color = 2'b11;
      12'hbb7: color = 2'b11;
      12'hbb8: color = 2'b11;
      12'hbb9: color = 2'b11;
      12'hbba: color = 2'b11;
      12'hbbb: color = 2'b00;
      12'hbbc: color = 2'b00;
      12'hbbd: color = 2'b00;
      12'hbbe: color = 2'b11;
      12'hbbf: color = 2'b11;
      12'hbc0: color = 2'b11;
      12'hbc1: color = 2'b11;
      12'hbc2: color = 2'b00;
      12'hbc3: color = 2'b00;
      12'hbc4: color = 2'b00;
      12'hbc5: color = 2'b00;
      12'hbc6: color = 2'b00;
      12'hbc7: color = 2'b00;
      12'hbc8: color = 2'b00;
      12'hbc9: color = 2'b11;
      12'hbca: color = 2'b11;
      12'hbcb: color = 2'b11;
      12'hbcc: color = 2'b11;
      12'hbcd: color = 2'b11;
      12'hbce: color = 2'b00;
      12'hbcf: color = 2'b00;
      12'hbd0: color = 2'b01;
      12'hbd1: color = 2'b01;
      12'hbd2: color = 2'b01;
      12'hbd3: color = 2'b01;
      12'hbd4: color = 2'b01;
      12'hbd5: color = 2'b01;
      12'hbd6: color = 2'b01;
      12'hbd7: color = 2'b00;
      12'hbd8: color = 2'b00;
      12'hbd9: color = 2'b01;
      12'hbda: color = 2'b01;
      12'hbdb: color = 2'b01;
      12'hbdc: color = 2'b01;
      12'hbdd: color = 2'b01;
      12'hbde: color = 2'b01;
      12'hbdf: color = 2'b01;
      12'hbe0: color = 2'b00;
      12'hbe1: color = 2'b00;
      12'hbe2: color = 2'b10;
      12'hbe3: color = 2'b10;
      12'hbe4: color = 2'b10;
      12'hbe5: color = 2'b10;
      12'hbe6: color = 2'b10;
      12'hbe7: color = 2'b00;
      12'hbe8: color = 2'b00;
      12'hbe9: color = 2'b11;
      12'hbea: color = 2'b11;
      12'hbeb: color = 2'b11;
      12'hbec: color = 2'b11;
      12'hbed: color = 2'b11;
      12'hbee: color = 2'b11;
      12'hbef: color = 2'b11;
      12'hbf0: color = 2'b00;
      12'hbf1: color = 2'b00;
      12'hbf2: color = 2'b00;
      12'hbf3: color = 2'b00;
      12'hbf4: color = 2'b00;
      12'hbf5: color = 2'b11;
      12'hbf6: color = 2'b11;
      12'hbf7: color = 2'b11;
      12'hbf8: color = 2'b11;
      12'hbf9: color = 2'b11;
      12'hbfa: color = 2'b11;
      12'hbfb: color = 2'b00;
      12'hbfc: color = 2'b00;
      12'hbfd: color = 2'b00;
      12'hbfe: color = 2'b11;
      12'hbff: color = 2'b11;
      12'hc00: color = 2'b00;
      12'hc01: color = 2'b00;
      12'hc02: color = 2'b11;
      12'hc03: color = 2'b11;
      12'hc04: color = 2'b11;
      12'hc05: color = 2'b01;
      12'hc06: color = 2'b01;
      12'hc07: color = 2'b01;
      12'hc08: color = 2'b01;
      12'hc09: color = 2'b00;
      12'hc0a: color = 2'b00;
      12'hc0b: color = 2'b00;
      12'hc0c: color = 2'b00;
      12'hc0d: color = 2'b00;
      12'hc0e: color = 2'b00;
      12'hc0f: color = 2'b00;
      12'hc10: color = 2'b00;
      12'hc11: color = 2'b00;
      12'hc12: color = 2'b00;
      12'hc13: color = 2'b00;
      12'hc14: color = 2'b00;
      12'hc15: color = 2'b00;
      12'hc16: color = 2'b00;
      12'hc17: color = 2'b01;
      12'hc18: color = 2'b01;
      12'hc19: color = 2'b01;
      12'hc1a: color = 2'b01;
      12'hc1b: color = 2'b01;
      12'hc1c: color = 2'b01;
      12'hc1d: color = 2'b01;
      12'hc1e: color = 2'b01;
      12'hc1f: color = 2'b01;
      12'hc20: color = 2'b00;
      12'hc21: color = 2'b00;
      12'hc22: color = 2'b10;
      12'hc23: color = 2'b10;
      12'hc24: color = 2'b10;
      12'hc25: color = 2'b00;
      12'hc26: color = 2'b00;
      12'hc27: color = 2'b10;
      12'hc28: color = 2'b10;
      12'hc29: color = 2'b11;
      12'hc2a: color = 2'b11;
      12'hc2b: color = 2'b11;
      12'hc2c: color = 2'b11;
      12'hc2d: color = 2'b11;
      12'hc2e: color = 2'b11;
      12'hc2f: color = 2'b11;
      12'hc30: color = 2'b00;
      12'hc31: color = 2'b00;
      12'hc32: color = 2'b10;
      12'hc33: color = 2'b10;
      12'hc34: color = 2'b10;
      12'hc35: color = 2'b11;
      12'hc36: color = 2'b11;
      12'hc37: color = 2'b11;
      12'hc38: color = 2'b11;
      12'hc39: color = 2'b11;
      12'hc3a: color = 2'b11;
      12'hc3b: color = 2'b00;
      12'hc3c: color = 2'b00;
      12'hc3d: color = 2'b00;
      12'hc3e: color = 2'b11;
      12'hc3f: color = 2'b11;
      12'hc40: color = 2'b00;
      12'hc41: color = 2'b00;
      12'hc42: color = 2'b11;
      12'hc43: color = 2'b11;
      12'hc44: color = 2'b11;
      12'hc45: color = 2'b01;
      12'hc46: color = 2'b01;
      12'hc47: color = 2'b01;
      12'hc48: color = 2'b01;
      12'hc49: color = 2'b00;
      12'hc4a: color = 2'b00;
      12'hc4b: color = 2'b00;
      12'hc4c: color = 2'b00;
      12'hc4d: color = 2'b00;
      12'hc4e: color = 2'b00;
      12'hc4f: color = 2'b00;
      12'hc50: color = 2'b00;
      12'hc51: color = 2'b00;
      12'hc52: color = 2'b00;
      12'hc53: color = 2'b00;
      12'hc54: color = 2'b00;
      12'hc55: color = 2'b00;
      12'hc56: color = 2'b00;
      12'hc57: color = 2'b01;
      12'hc58: color = 2'b01;
      12'hc59: color = 2'b01;
      12'hc5a: color = 2'b01;
      12'hc5b: color = 2'b01;
      12'hc5c: color = 2'b01;
      12'hc5d: color = 2'b01;
      12'hc5e: color = 2'b01;
      12'hc5f: color = 2'b01;
      12'hc60: color = 2'b00;
      12'hc61: color = 2'b00;
      12'hc62: color = 2'b10;
      12'hc63: color = 2'b10;
      12'hc64: color = 2'b10;
      12'hc65: color = 2'b00;
      12'hc66: color = 2'b00;
      12'hc67: color = 2'b10;
      12'hc68: color = 2'b10;
      12'hc69: color = 2'b11;
      12'hc6a: color = 2'b11;
      12'hc6b: color = 2'b11;
      12'hc6c: color = 2'b11;
      12'hc6d: color = 2'b11;
      12'hc6e: color = 2'b11;
      12'hc6f: color = 2'b11;
      12'hc70: color = 2'b00;
      12'hc71: color = 2'b00;
      12'hc72: color = 2'b10;
      12'hc73: color = 2'b10;
      12'hc74: color = 2'b10;
      12'hc75: color = 2'b11;
      12'hc76: color = 2'b11;
      12'hc77: color = 2'b11;
      12'hc78: color = 2'b11;
      12'hc79: color = 2'b11;
      12'hc7a: color = 2'b11;
      12'hc7b: color = 2'b00;
      12'hc7c: color = 2'b00;
      12'hc7d: color = 2'b00;
      12'hc7e: color = 2'b11;
      12'hc7f: color = 2'b11;
      12'hc80: color = 2'b00;
      12'hc81: color = 2'b00;
      12'hc82: color = 2'b00;
      12'hc83: color = 2'b00;
      12'hc84: color = 2'b00;
      12'hc85: color = 2'b01;
      12'hc86: color = 2'b01;
      12'hc87: color = 2'b01;
      12'hc88: color = 2'b01;
      12'hc89: color = 2'b01;
      12'hc8a: color = 2'b01;
      12'hc8b: color = 2'b01;
      12'hc8c: color = 2'b01;
      12'hc8d: color = 2'b01;
      12'hc8e: color = 2'b01;
      12'hc8f: color = 2'b01;
      12'hc90: color = 2'b01;
      12'hc91: color = 2'b01;
      12'hc92: color = 2'b00;
      12'hc93: color = 2'b00;
      12'hc94: color = 2'b00;
      12'hc95: color = 2'b00;
      12'hc96: color = 2'b00;
      12'hc97: color = 2'b01;
      12'hc98: color = 2'b01;
      12'hc99: color = 2'b01;
      12'hc9a: color = 2'b01;
      12'hc9b: color = 2'b01;
      12'hc9c: color = 2'b01;
      12'hc9d: color = 2'b01;
      12'hc9e: color = 2'b00;
      12'hc9f: color = 2'b00;
      12'hca0: color = 2'b10;
      12'hca1: color = 2'b10;
      12'hca2: color = 2'b10;
      12'hca3: color = 2'b10;
      12'hca4: color = 2'b10;
      12'hca5: color = 2'b00;
      12'hca6: color = 2'b00;
      12'hca7: color = 2'b10;
      12'hca8: color = 2'b10;
      12'hca9: color = 2'b10;
      12'hcaa: color = 2'b10;
      12'hcab: color = 2'b11;
      12'hcac: color = 2'b11;
      12'hcad: color = 2'b11;
      12'hcae: color = 2'b11;
      12'hcaf: color = 2'b11;
      12'hcb0: color = 2'b11;
      12'hcb1: color = 2'b11;
      12'hcb2: color = 2'b01;
      12'hcb3: color = 2'b01;
      12'hcb4: color = 2'b01;
      12'hcb5: color = 2'b01;
      12'hcb6: color = 2'b01;
      12'hcb7: color = 2'b11;
      12'hcb8: color = 2'b11;
      12'hcb9: color = 2'b11;
      12'hcba: color = 2'b11;
      12'hcbb: color = 2'b11;
      12'hcbc: color = 2'b11;
      12'hcbd: color = 2'b11;
      12'hcbe: color = 2'b01;
      12'hcbf: color = 2'b01;
      12'hcc0: color = 2'b00;
      12'hcc1: color = 2'b00;
      12'hcc2: color = 2'b00;
      12'hcc3: color = 2'b00;
      12'hcc4: color = 2'b00;
      12'hcc5: color = 2'b01;
      12'hcc6: color = 2'b01;
      12'hcc7: color = 2'b01;
      12'hcc8: color = 2'b01;
      12'hcc9: color = 2'b01;
      12'hcca: color = 2'b01;
      12'hccb: color = 2'b01;
      12'hccc: color = 2'b01;
      12'hccd: color = 2'b01;
      12'hcce: color = 2'b01;
      12'hccf: color = 2'b01;
      12'hcd0: color = 2'b01;
      12'hcd1: color = 2'b01;
      12'hcd2: color = 2'b00;
      12'hcd3: color = 2'b00;
      12'hcd4: color = 2'b00;
      12'hcd5: color = 2'b00;
      12'hcd6: color = 2'b00;
      12'hcd7: color = 2'b01;
      12'hcd8: color = 2'b01;
      12'hcd9: color = 2'b01;
      12'hcda: color = 2'b01;
      12'hcdb: color = 2'b01;
      12'hcdc: color = 2'b01;
      12'hcdd: color = 2'b01;
      12'hcde: color = 2'b00;
      12'hcdf: color = 2'b00;
      12'hce0: color = 2'b10;
      12'hce1: color = 2'b10;
      12'hce2: color = 2'b10;
      12'hce3: color = 2'b10;
      12'hce4: color = 2'b10;
      12'hce5: color = 2'b00;
      12'hce6: color = 2'b00;
      12'hce7: color = 2'b10;
      12'hce8: color = 2'b10;
      12'hce9: color = 2'b10;
      12'hcea: color = 2'b10;
      12'hceb: color = 2'b11;
      12'hcec: color = 2'b11;
      12'hced: color = 2'b11;
      12'hcee: color = 2'b11;
      12'hcef: color = 2'b11;
      12'hcf0: color = 2'b11;
      12'hcf1: color = 2'b11;
      12'hcf2: color = 2'b01;
      12'hcf3: color = 2'b01;
      12'hcf4: color = 2'b01;
      12'hcf5: color = 2'b01;
      12'hcf6: color = 2'b01;
      12'hcf7: color = 2'b11;
      12'hcf8: color = 2'b11;
      12'hcf9: color = 2'b11;
      12'hcfa: color = 2'b11;
      12'hcfb: color = 2'b11;
      12'hcfc: color = 2'b11;
      12'hcfd: color = 2'b11;
      12'hcfe: color = 2'b01;
      12'hcff: color = 2'b01;
      12'hd00: color = 2'b00;
      12'hd01: color = 2'b00;
      12'hd02: color = 2'b00;
      12'hd03: color = 2'b00;
      12'hd04: color = 2'b00;
      12'hd05: color = 2'b01;
      12'hd06: color = 2'b01;
      12'hd07: color = 2'b01;
      12'hd08: color = 2'b01;
      12'hd09: color = 2'b01;
      12'hd0a: color = 2'b01;
      12'hd0b: color = 2'b01;
      12'hd0c: color = 2'b01;
      12'hd0d: color = 2'b01;
      12'hd0e: color = 2'b01;
      12'hd0f: color = 2'b01;
      12'hd10: color = 2'b01;
      12'hd11: color = 2'b01;
      12'hd12: color = 2'b01;
      12'hd13: color = 2'b01;
      12'hd14: color = 2'b01;
      12'hd15: color = 2'b00;
      12'hd16: color = 2'b00;
      12'hd17: color = 2'b01;
      12'hd18: color = 2'b01;
      12'hd19: color = 2'b01;
      12'hd1a: color = 2'b01;
      12'hd1b: color = 2'b01;
      12'hd1c: color = 2'b01;
      12'hd1d: color = 2'b01;
      12'hd1e: color = 2'b00;
      12'hd1f: color = 2'b00;
      12'hd20: color = 2'b00;
      12'hd21: color = 2'b00;
      12'hd22: color = 2'b00;
      12'hd23: color = 2'b00;
      12'hd24: color = 2'b00;
      12'hd25: color = 2'b10;
      12'hd26: color = 2'b10;
      12'hd27: color = 2'b10;
      12'hd28: color = 2'b10;
      12'hd29: color = 2'b10;
      12'hd2a: color = 2'b10;
      12'hd2b: color = 2'b10;
      12'hd2c: color = 2'b10;
      12'hd2d: color = 2'b10;
      12'hd2e: color = 2'b11;
      12'hd2f: color = 2'b11;
      12'hd30: color = 2'b11;
      12'hd31: color = 2'b11;
      12'hd32: color = 2'b00;
      12'hd33: color = 2'b00;
      12'hd34: color = 2'b00;
      12'hd35: color = 2'b11;
      12'hd36: color = 2'b11;
      12'hd37: color = 2'b01;
      12'hd38: color = 2'b01;
      12'hd39: color = 2'b11;
      12'hd3a: color = 2'b11;
      12'hd3b: color = 2'b11;
      12'hd3c: color = 2'b11;
      12'hd3d: color = 2'b11;
      12'hd3e: color = 2'b00;
      12'hd3f: color = 2'b00;
      12'hd40: color = 2'b00;
      12'hd41: color = 2'b00;
      12'hd42: color = 2'b00;
      12'hd43: color = 2'b00;
      12'hd44: color = 2'b00;
      12'hd45: color = 2'b01;
      12'hd46: color = 2'b01;
      12'hd47: color = 2'b01;
      12'hd48: color = 2'b01;
      12'hd49: color = 2'b01;
      12'hd4a: color = 2'b01;
      12'hd4b: color = 2'b01;
      12'hd4c: color = 2'b01;
      12'hd4d: color = 2'b01;
      12'hd4e: color = 2'b01;
      12'hd4f: color = 2'b01;
      12'hd50: color = 2'b01;
      12'hd51: color = 2'b01;
      12'hd52: color = 2'b01;
      12'hd53: color = 2'b01;
      12'hd54: color = 2'b01;
      12'hd55: color = 2'b00;
      12'hd56: color = 2'b00;
      12'hd57: color = 2'b01;
      12'hd58: color = 2'b01;
      12'hd59: color = 2'b01;
      12'hd5a: color = 2'b01;
      12'hd5b: color = 2'b01;
      12'hd5c: color = 2'b01;
      12'hd5d: color = 2'b01;
      12'hd5e: color = 2'b00;
      12'hd5f: color = 2'b00;
      12'hd60: color = 2'b00;
      12'hd61: color = 2'b00;
      12'hd62: color = 2'b00;
      12'hd63: color = 2'b00;
      12'hd64: color = 2'b00;
      12'hd65: color = 2'b10;
      12'hd66: color = 2'b10;
      12'hd67: color = 2'b10;
      12'hd68: color = 2'b10;
      12'hd69: color = 2'b10;
      12'hd6a: color = 2'b10;
      12'hd6b: color = 2'b10;
      12'hd6c: color = 2'b10;
      12'hd6d: color = 2'b10;
      12'hd6e: color = 2'b11;
      12'hd6f: color = 2'b11;
      12'hd70: color = 2'b11;
      12'hd71: color = 2'b11;
      12'hd72: color = 2'b00;
      12'hd73: color = 2'b00;
      12'hd74: color = 2'b00;
      12'hd75: color = 2'b11;
      12'hd76: color = 2'b11;
      12'hd77: color = 2'b01;
      12'hd78: color = 2'b01;
      12'hd79: color = 2'b11;
      12'hd7a: color = 2'b11;
      12'hd7b: color = 2'b11;
      12'hd7c: color = 2'b11;
      12'hd7d: color = 2'b11;
      12'hd7e: color = 2'b00;
      12'hd7f: color = 2'b00;
      12'hd80: color = 2'b00;
      12'hd81: color = 2'b00;
      12'hd82: color = 2'b00;
      12'hd83: color = 2'b00;
      12'hd84: color = 2'b00;
      12'hd85: color = 2'b01;
      12'hd86: color = 2'b01;
      12'hd87: color = 2'b01;
      12'hd88: color = 2'b01;
      12'hd89: color = 2'b01;
      12'hd8a: color = 2'b01;
      12'hd8b: color = 2'b01;
      12'hd8c: color = 2'b01;
      12'hd8d: color = 2'b01;
      12'hd8e: color = 2'b01;
      12'hd8f: color = 2'b01;
      12'hd90: color = 2'b01;
      12'hd91: color = 2'b01;
      12'hd92: color = 2'b01;
      12'hd93: color = 2'b01;
      12'hd94: color = 2'b01;
      12'hd95: color = 2'b00;
      12'hd96: color = 2'b00;
      12'hd97: color = 2'b01;
      12'hd98: color = 2'b01;
      12'hd99: color = 2'b01;
      12'hd9a: color = 2'b01;
      12'hd9b: color = 2'b01;
      12'hd9c: color = 2'b01;
      12'hd9d: color = 2'b01;
      12'hd9e: color = 2'b00;
      12'hd9f: color = 2'b00;
      12'hda0: color = 2'b00;
      12'hda1: color = 2'b00;
      12'hda2: color = 2'b00;
      12'hda3: color = 2'b00;
      12'hda4: color = 2'b00;
      12'hda5: color = 2'b10;
      12'hda6: color = 2'b10;
      12'hda7: color = 2'b10;
      12'hda8: color = 2'b10;
      12'hda9: color = 2'b10;
      12'hdaa: color = 2'b10;
      12'hdab: color = 2'b10;
      12'hdac: color = 2'b10;
      12'hdad: color = 2'b10;
      12'hdae: color = 2'b11;
      12'hdaf: color = 2'b11;
      12'hdb0: color = 2'b11;
      12'hdb1: color = 2'b11;
      12'hdb2: color = 2'b00;
      12'hdb3: color = 2'b00;
      12'hdb4: color = 2'b00;
      12'hdb5: color = 2'b11;
      12'hdb6: color = 2'b11;
      12'hdb7: color = 2'b01;
      12'hdb8: color = 2'b01;
      12'hdb9: color = 2'b11;
      12'hdba: color = 2'b11;
      12'hdbb: color = 2'b11;
      12'hdbc: color = 2'b11;
      12'hdbd: color = 2'b11;
      12'hdbe: color = 2'b00;
      12'hdbf: color = 2'b00;
      12'hdc0: color = 2'b11;
      12'hdc1: color = 2'b11;
      12'hdc2: color = 2'b00;
      12'hdc3: color = 2'b00;
      12'hdc4: color = 2'b00;
      12'hdc5: color = 2'b01;
      12'hdc6: color = 2'b01;
      12'hdc7: color = 2'b01;
      12'hdc8: color = 2'b01;
      12'hdc9: color = 2'b01;
      12'hdca: color = 2'b01;
      12'hdcb: color = 2'b01;
      12'hdcc: color = 2'b01;
      12'hdcd: color = 2'b01;
      12'hdce: color = 2'b01;
      12'hdcf: color = 2'b01;
      12'hdd0: color = 2'b01;
      12'hdd1: color = 2'b01;
      12'hdd2: color = 2'b01;
      12'hdd3: color = 2'b01;
      12'hdd4: color = 2'b01;
      12'hdd5: color = 2'b00;
      12'hdd6: color = 2'b00;
      12'hdd7: color = 2'b01;
      12'hdd8: color = 2'b01;
      12'hdd9: color = 2'b01;
      12'hdda: color = 2'b01;
      12'hddb: color = 2'b00;
      12'hddc: color = 2'b00;
      12'hddd: color = 2'b00;
      12'hdde: color = 2'b01;
      12'hddf: color = 2'b01;
      12'hde0: color = 2'b01;
      12'hde1: color = 2'b01;
      12'hde2: color = 2'b00;
      12'hde3: color = 2'b00;
      12'hde4: color = 2'b00;
      12'hde5: color = 2'b10;
      12'hde6: color = 2'b10;
      12'hde7: color = 2'b10;
      12'hde8: color = 2'b10;
      12'hde9: color = 2'b10;
      12'hdea: color = 2'b10;
      12'hdeb: color = 2'b10;
      12'hdec: color = 2'b10;
      12'hded: color = 2'b10;
      12'hdee: color = 2'b10;
      12'hdef: color = 2'b10;
      12'hdf0: color = 2'b10;
      12'hdf1: color = 2'b10;
      12'hdf2: color = 2'b00;
      12'hdf3: color = 2'b00;
      12'hdf4: color = 2'b00;
      12'hdf5: color = 2'b11;
      12'hdf6: color = 2'b11;
      12'hdf7: color = 2'b11;
      12'hdf8: color = 2'b11;
      12'hdf9: color = 2'b00;
      12'hdfa: color = 2'b00;
      12'hdfb: color = 2'b10;
      12'hdfc: color = 2'b10;
      12'hdfd: color = 2'b10;
      12'hdfe: color = 2'b00;
      12'hdff: color = 2'b00;
      12'he00: color = 2'b11;
      12'he01: color = 2'b11;
      12'he02: color = 2'b00;
      12'he03: color = 2'b00;
      12'he04: color = 2'b00;
      12'he05: color = 2'b01;
      12'he06: color = 2'b01;
      12'he07: color = 2'b01;
      12'he08: color = 2'b01;
      12'he09: color = 2'b01;
      12'he0a: color = 2'b01;
      12'he0b: color = 2'b01;
      12'he0c: color = 2'b01;
      12'he0d: color = 2'b01;
      12'he0e: color = 2'b01;
      12'he0f: color = 2'b01;
      12'he10: color = 2'b01;
      12'he11: color = 2'b01;
      12'he12: color = 2'b01;
      12'he13: color = 2'b01;
      12'he14: color = 2'b01;
      12'he15: color = 2'b00;
      12'he16: color = 2'b00;
      12'he17: color = 2'b01;
      12'he18: color = 2'b01;
      12'he19: color = 2'b01;
      12'he1a: color = 2'b01;
      12'he1b: color = 2'b00;
      12'he1c: color = 2'b00;
      12'he1d: color = 2'b00;
      12'he1e: color = 2'b01;
      12'he1f: color = 2'b01;
      12'he20: color = 2'b01;
      12'he21: color = 2'b01;
      12'he22: color = 2'b00;
      12'he23: color = 2'b00;
      12'he24: color = 2'b00;
      12'he25: color = 2'b10;
      12'he26: color = 2'b10;
      12'he27: color = 2'b10;
      12'he28: color = 2'b10;
      12'he29: color = 2'b10;
      12'he2a: color = 2'b10;
      12'he2b: color = 2'b10;
      12'he2c: color = 2'b10;
      12'he2d: color = 2'b10;
      12'he2e: color = 2'b10;
      12'he2f: color = 2'b10;
      12'he30: color = 2'b10;
      12'he31: color = 2'b10;
      12'he32: color = 2'b00;
      12'he33: color = 2'b00;
      12'he34: color = 2'b00;
      12'he35: color = 2'b11;
      12'he36: color = 2'b11;
      12'he37: color = 2'b11;
      12'he38: color = 2'b11;
      12'he39: color = 2'b00;
      12'he3a: color = 2'b00;
      12'he3b: color = 2'b10;
      12'he3c: color = 2'b10;
      12'he3d: color = 2'b10;
      12'he3e: color = 2'b00;
      12'he3f: color = 2'b00;
      12'he40: color = 2'b11;
      12'he41: color = 2'b11;
      12'he42: color = 2'b00;
      12'he43: color = 2'b00;
      12'he44: color = 2'b00;
      12'he45: color = 2'b01;
      12'he46: color = 2'b01;
      12'he47: color = 2'b01;
      12'he48: color = 2'b01;
      12'he49: color = 2'b01;
      12'he4a: color = 2'b01;
      12'he4b: color = 2'b01;
      12'he4c: color = 2'b01;
      12'he4d: color = 2'b01;
      12'he4e: color = 2'b01;
      12'he4f: color = 2'b01;
      12'he50: color = 2'b01;
      12'he51: color = 2'b01;
      12'he52: color = 2'b01;
      12'he53: color = 2'b01;
      12'he54: color = 2'b01;
      12'he55: color = 2'b00;
      12'he56: color = 2'b00;
      12'he57: color = 2'b01;
      12'he58: color = 2'b01;
      12'he59: color = 2'b01;
      12'he5a: color = 2'b01;
      12'he5b: color = 2'b00;
      12'he5c: color = 2'b00;
      12'he5d: color = 2'b00;
      12'he5e: color = 2'b01;
      12'he5f: color = 2'b01;
      12'he60: color = 2'b00;
      12'he61: color = 2'b00;
      12'he62: color = 2'b10;
      12'he63: color = 2'b10;
      12'he64: color = 2'b10;
      12'he65: color = 2'b00;
      12'he66: color = 2'b00;
      12'he67: color = 2'b10;
      12'he68: color = 2'b10;
      12'he69: color = 2'b10;
      12'he6a: color = 2'b10;
      12'he6b: color = 2'b10;
      12'he6c: color = 2'b10;
      12'he6d: color = 2'b10;
      12'he6e: color = 2'b10;
      12'he6f: color = 2'b10;
      12'he70: color = 2'b10;
      12'he71: color = 2'b10;
      12'he72: color = 2'b00;
      12'he73: color = 2'b00;
      12'he74: color = 2'b00;
      12'he75: color = 2'b11;
      12'he76: color = 2'b11;
      12'he77: color = 2'b00;
      12'he78: color = 2'b00;
      12'he79: color = 2'b00;
      12'he7a: color = 2'b00;
      12'he7b: color = 2'b00;
      12'he7c: color = 2'b00;
      12'he7d: color = 2'b00;
      12'he7e: color = 2'b11;
      12'he7f: color = 2'b11;
      12'he80: color = 2'b11;
      12'he81: color = 2'b11;
      12'he82: color = 2'b00;
      12'he83: color = 2'b00;
      12'he84: color = 2'b00;
      12'he85: color = 2'b01;
      12'he86: color = 2'b01;
      12'he87: color = 2'b01;
      12'he88: color = 2'b01;
      12'he89: color = 2'b01;
      12'he8a: color = 2'b01;
      12'he8b: color = 2'b01;
      12'he8c: color = 2'b01;
      12'he8d: color = 2'b01;
      12'he8e: color = 2'b01;
      12'he8f: color = 2'b01;
      12'he90: color = 2'b01;
      12'he91: color = 2'b01;
      12'he92: color = 2'b01;
      12'he93: color = 2'b01;
      12'he94: color = 2'b01;
      12'he95: color = 2'b00;
      12'he96: color = 2'b00;
      12'he97: color = 2'b01;
      12'he98: color = 2'b01;
      12'he99: color = 2'b01;
      12'he9a: color = 2'b01;
      12'he9b: color = 2'b00;
      12'he9c: color = 2'b00;
      12'he9d: color = 2'b00;
      12'he9e: color = 2'b01;
      12'he9f: color = 2'b01;
      12'hea0: color = 2'b00;
      12'hea1: color = 2'b00;
      12'hea2: color = 2'b10;
      12'hea3: color = 2'b10;
      12'hea4: color = 2'b10;
      12'hea5: color = 2'b00;
      12'hea6: color = 2'b00;
      12'hea7: color = 2'b10;
      12'hea8: color = 2'b10;
      12'hea9: color = 2'b10;
      12'heaa: color = 2'b10;
      12'heab: color = 2'b10;
      12'heac: color = 2'b10;
      12'head: color = 2'b10;
      12'heae: color = 2'b10;
      12'heaf: color = 2'b10;
      12'heb0: color = 2'b10;
      12'heb1: color = 2'b10;
      12'heb2: color = 2'b00;
      12'heb3: color = 2'b00;
      12'heb4: color = 2'b00;
      12'heb5: color = 2'b11;
      12'heb6: color = 2'b11;
      12'heb7: color = 2'b00;
      12'heb8: color = 2'b00;
      12'heb9: color = 2'b00;
      12'heba: color = 2'b00;
      12'hebb: color = 2'b00;
      12'hebc: color = 2'b00;
      12'hebd: color = 2'b00;
      12'hebe: color = 2'b11;
      12'hebf: color = 2'b11;
      12'hec0: color = 2'b11;
      12'hec1: color = 2'b11;
      12'hec2: color = 2'b11;
      12'hec3: color = 2'b11;
      12'hec4: color = 2'b11;
      12'hec5: color = 2'b00;
      12'hec6: color = 2'b00;
      12'hec7: color = 2'b00;
      12'hec8: color = 2'b00;
      12'hec9: color = 2'b01;
      12'heca: color = 2'b01;
      12'hecb: color = 2'b01;
      12'hecc: color = 2'b01;
      12'hecd: color = 2'b01;
      12'hece: color = 2'b01;
      12'hecf: color = 2'b01;
      12'hed0: color = 2'b01;
      12'hed1: color = 2'b01;
      12'hed2: color = 2'b01;
      12'hed3: color = 2'b01;
      12'hed4: color = 2'b01;
      12'hed5: color = 2'b01;
      12'hed6: color = 2'b01;
      12'hed7: color = 2'b00;
      12'hed8: color = 2'b00;
      12'hed9: color = 2'b00;
      12'heda: color = 2'b00;
      12'hedb: color = 2'b01;
      12'hedc: color = 2'b01;
      12'hedd: color = 2'b01;
      12'hede: color = 2'b00;
      12'hedf: color = 2'b00;
      12'hee0: color = 2'b10;
      12'hee1: color = 2'b10;
      12'hee2: color = 2'b00;
      12'hee3: color = 2'b00;
      12'hee4: color = 2'b00;
      12'hee5: color = 2'b11;
      12'hee6: color = 2'b11;
      12'hee7: color = 2'b00;
      12'hee8: color = 2'b00;
      12'hee9: color = 2'b10;
      12'heea: color = 2'b10;
      12'heeb: color = 2'b10;
      12'heec: color = 2'b10;
      12'heed: color = 2'b10;
      12'heee: color = 2'b10;
      12'heef: color = 2'b10;
      12'hef0: color = 2'b00;
      12'hef1: color = 2'b00;
      12'hef2: color = 2'b00;
      12'hef3: color = 2'b00;
      12'hef4: color = 2'b00;
      12'hef5: color = 2'b00;
      12'hef6: color = 2'b00;
      12'hef7: color = 2'b11;
      12'hef8: color = 2'b11;
      12'hef9: color = 2'b11;
      12'hefa: color = 2'b11;
      12'hefb: color = 2'b11;
      12'hefc: color = 2'b11;
      12'hefd: color = 2'b11;
      12'hefe: color = 2'b11;
      12'heff: color = 2'b11;
      12'hf00: color = 2'b11;
      12'hf01: color = 2'b11;
      12'hf02: color = 2'b11;
      12'hf03: color = 2'b11;
      12'hf04: color = 2'b11;
      12'hf05: color = 2'b00;
      12'hf06: color = 2'b00;
      12'hf07: color = 2'b00;
      12'hf08: color = 2'b00;
      12'hf09: color = 2'b01;
      12'hf0a: color = 2'b01;
      12'hf0b: color = 2'b01;
      12'hf0c: color = 2'b01;
      12'hf0d: color = 2'b01;
      12'hf0e: color = 2'b01;
      12'hf0f: color = 2'b01;
      12'hf10: color = 2'b01;
      12'hf11: color = 2'b01;
      12'hf12: color = 2'b01;
      12'hf13: color = 2'b01;
      12'hf14: color = 2'b01;
      12'hf15: color = 2'b01;
      12'hf16: color = 2'b01;
      12'hf17: color = 2'b00;
      12'hf18: color = 2'b00;
      12'hf19: color = 2'b00;
      12'hf1a: color = 2'b00;
      12'hf1b: color = 2'b01;
      12'hf1c: color = 2'b01;
      12'hf1d: color = 2'b01;
      12'hf1e: color = 2'b00;
      12'hf1f: color = 2'b00;
      12'hf20: color = 2'b10;
      12'hf21: color = 2'b10;
      12'hf22: color = 2'b00;
      12'hf23: color = 2'b00;
      12'hf24: color = 2'b00;
      12'hf25: color = 2'b11;
      12'hf26: color = 2'b11;
      12'hf27: color = 2'b00;
      12'hf28: color = 2'b00;
      12'hf29: color = 2'b10;
      12'hf2a: color = 2'b10;
      12'hf2b: color = 2'b10;
      12'hf2c: color = 2'b10;
      12'hf2d: color = 2'b10;
      12'hf2e: color = 2'b10;
      12'hf2f: color = 2'b10;
      12'hf30: color = 2'b00;
      12'hf31: color = 2'b00;
      12'hf32: color = 2'b00;
      12'hf33: color = 2'b00;
      12'hf34: color = 2'b00;
      12'hf35: color = 2'b00;
      12'hf36: color = 2'b00;
      12'hf37: color = 2'b11;
      12'hf38: color = 2'b11;
      12'hf39: color = 2'b11;
      12'hf3a: color = 2'b11;
      12'hf3b: color = 2'b11;
      12'hf3c: color = 2'b11;
      12'hf3d: color = 2'b11;
      12'hf3e: color = 2'b11;
      12'hf3f: color = 2'b11;
      12'hf40: color = 2'b11;
      12'hf41: color = 2'b11;
      12'hf42: color = 2'b11;
      12'hf43: color = 2'b11;
      12'hf44: color = 2'b11;
      12'hf45: color = 2'b00;
      12'hf46: color = 2'b00;
      12'hf47: color = 2'b00;
      12'hf48: color = 2'b00;
      12'hf49: color = 2'b01;
      12'hf4a: color = 2'b01;
      12'hf4b: color = 2'b01;
      12'hf4c: color = 2'b01;
      12'hf4d: color = 2'b01;
      12'hf4e: color = 2'b01;
      12'hf4f: color = 2'b01;
      12'hf50: color = 2'b01;
      12'hf51: color = 2'b01;
      12'hf52: color = 2'b01;
      12'hf53: color = 2'b01;
      12'hf54: color = 2'b01;
      12'hf55: color = 2'b01;
      12'hf56: color = 2'b01;
      12'hf57: color = 2'b00;
      12'hf58: color = 2'b00;
      12'hf59: color = 2'b00;
      12'hf5a: color = 2'b00;
      12'hf5b: color = 2'b01;
      12'hf5c: color = 2'b01;
      12'hf5d: color = 2'b01;
      12'hf5e: color = 2'b00;
      12'hf5f: color = 2'b00;
      12'hf60: color = 2'b10;
      12'hf61: color = 2'b10;
      12'hf62: color = 2'b00;
      12'hf63: color = 2'b00;
      12'hf64: color = 2'b00;
      12'hf65: color = 2'b11;
      12'hf66: color = 2'b11;
      12'hf67: color = 2'b00;
      12'hf68: color = 2'b00;
      12'hf69: color = 2'b10;
      12'hf6a: color = 2'b10;
      12'hf6b: color = 2'b10;
      12'hf6c: color = 2'b10;
      12'hf6d: color = 2'b10;
      12'hf6e: color = 2'b10;
      12'hf6f: color = 2'b10;
      12'hf70: color = 2'b00;
      12'hf71: color = 2'b00;
      12'hf72: color = 2'b00;
      12'hf73: color = 2'b00;
      12'hf74: color = 2'b00;
      12'hf75: color = 2'b00;
      12'hf76: color = 2'b00;
      12'hf77: color = 2'b11;
      12'hf78: color = 2'b11;
      12'hf79: color = 2'b11;
      12'hf7a: color = 2'b11;
      12'hf7b: color = 2'b11;
      12'hf7c: color = 2'b11;
      12'hf7d: color = 2'b11;
      12'hf7e: color = 2'b11;
      12'hf7f: color = 2'b11;
      12'hf80: color = 2'b11;
      12'hf81: color = 2'b11;
      12'hf82: color = 2'b11;
      12'hf83: color = 2'b11;
      12'hf84: color = 2'b11;
      12'hf85: color = 2'b11;
      12'hf86: color = 2'b11;
      12'hf87: color = 2'b11;
      12'hf88: color = 2'b11;
      12'hf89: color = 2'b00;
      12'hf8a: color = 2'b00;
      12'hf8b: color = 2'b00;
      12'hf8c: color = 2'b00;
      12'hf8d: color = 2'b00;
      12'hf8e: color = 2'b00;
      12'hf8f: color = 2'b00;
      12'hf90: color = 2'b00;
      12'hf91: color = 2'b00;
      12'hf92: color = 2'b00;
      12'hf93: color = 2'b00;
      12'hf94: color = 2'b00;
      12'hf95: color = 2'b00;
      12'hf96: color = 2'b00;
      12'hf97: color = 2'b01;
      12'hf98: color = 2'b01;
      12'hf99: color = 2'b00;
      12'hf9a: color = 2'b00;
      12'hf9b: color = 2'b01;
      12'hf9c: color = 2'b01;
      12'hf9d: color = 2'b01;
      12'hf9e: color = 2'b01;
      12'hf9f: color = 2'b01;
      12'hfa0: color = 2'b00;
      12'hfa1: color = 2'b00;
      12'hfa2: color = 2'b11;
      12'hfa3: color = 2'b11;
      12'hfa4: color = 2'b11;
      12'hfa5: color = 2'b11;
      12'hfa6: color = 2'b11;
      12'hfa7: color = 2'b11;
      12'hfa8: color = 2'b11;
      12'hfa9: color = 2'b00;
      12'hfaa: color = 2'b00;
      12'hfab: color = 2'b00;
      12'hfac: color = 2'b00;
      12'hfad: color = 2'b00;
      12'hfae: color = 2'b00;
      12'hfaf: color = 2'b00;
      12'hfb0: color = 2'b00;
      12'hfb1: color = 2'b00;
      12'hfb2: color = 2'b11;
      12'hfb3: color = 2'b11;
      12'hfb4: color = 2'b11;
      12'hfb5: color = 2'b11;
      12'hfb6: color = 2'b11;
      12'hfb7: color = 2'b11;
      12'hfb8: color = 2'b11;
      12'hfb9: color = 2'b11;
      12'hfba: color = 2'b11;
      12'hfbb: color = 2'b11;
      12'hfbc: color = 2'b11;
      12'hfbd: color = 2'b11;
      12'hfbe: color = 2'b11;
      12'hfbf: color = 2'b11;
      12'hfc0: color = 2'b11;
      12'hfc1: color = 2'b11;
      12'hfc2: color = 2'b11;
      12'hfc3: color = 2'b11;
      12'hfc4: color = 2'b11;
      12'hfc5: color = 2'b11;
      12'hfc6: color = 2'b11;
      12'hfc7: color = 2'b11;
      12'hfc8: color = 2'b11;
      12'hfc9: color = 2'b00;
      12'hfca: color = 2'b00;
      12'hfcb: color = 2'b00;
      12'hfcc: color = 2'b00;
      12'hfcd: color = 2'b00;
      12'hfce: color = 2'b00;
      12'hfcf: color = 2'b00;
      12'hfd0: color = 2'b00;
      12'hfd1: color = 2'b00;
      12'hfd2: color = 2'b00;
      12'hfd3: color = 2'b00;
      12'hfd4: color = 2'b00;
      12'hfd5: color = 2'b00;
      12'hfd6: color = 2'b00;
      12'hfd7: color = 2'b01;
      12'hfd8: color = 2'b01;
      12'hfd9: color = 2'b00;
      12'hfda: color = 2'b00;
      12'hfdb: color = 2'b01;
      12'hfdc: color = 2'b01;
      12'hfdd: color = 2'b01;
      12'hfde: color = 2'b01;
      12'hfdf: color = 2'b01;
      12'hfe0: color = 2'b00;
      12'hfe1: color = 2'b00;
      12'hfe2: color = 2'b11;
      12'hfe3: color = 2'b11;
      12'hfe4: color = 2'b11;
      12'hfe5: color = 2'b11;
      12'hfe6: color = 2'b11;
      12'hfe7: color = 2'b11;
      12'hfe8: color = 2'b11;
      12'hfe9: color = 2'b00;
      12'hfea: color = 2'b00;
      12'hfeb: color = 2'b00;
      12'hfec: color = 2'b00;
      12'hfed: color = 2'b00;
      12'hfee: color = 2'b00;
      12'hfef: color = 2'b00;
      12'hff0: color = 2'b00;
      12'hff1: color = 2'b00;
      12'hff2: color = 2'b11;
      12'hff3: color = 2'b11;
      12'hff4: color = 2'b11;
      12'hff5: color = 2'b11;
      12'hff6: color = 2'b11;
      12'hff7: color = 2'b11;
      12'hff8: color = 2'b11;
      12'hff9: color = 2'b11;
      12'hffa: color = 2'b11;
      12'hffb: color = 2'b11;
      12'hffc: color = 2'b11;
      12'hffd: color = 2'b11;
      12'hffe: color = 2'b11;
      12'hfff: color = 2'b11;
   endcase
end
endmodule
