module Desk
(
   input            clock, 
   input      [7:0] x,
   input      [7:0] y, 
   output reg [1:0] color
);

   reg [12:0] addr;
   always @( posedge clock )
      addr <= {y[5:0],x[6:0]};

always @(*) begin
   case( addr )
      13'h0000: color = 2'b11;
      13'h0001: color = 2'b11;
      13'h0002: color = 2'b11;
      13'h0003: color = 2'b11;
      13'h0004: color = 2'b10;
      13'h0005: color = 2'b10;
      13'h0006: color = 2'b11;
      13'h0007: color = 2'b11;
      13'h0008: color = 2'b10;
      13'h0009: color = 2'b10;
      13'h000a: color = 2'b11;
      13'h000b: color = 2'b11;
      13'h000c: color = 2'b11;
      13'h000d: color = 2'b11;
      13'h000e: color = 2'b11;
      13'h000f: color = 2'b11;
      13'h0010: color = 2'b11;
      13'h0011: color = 2'b11;
      13'h0012: color = 2'b11;
      13'h0013: color = 2'b11;
      13'h0014: color = 2'b10;
      13'h0015: color = 2'b10;
      13'h0016: color = 2'b11;
      13'h0017: color = 2'b11;
      13'h0018: color = 2'b10;
      13'h0019: color = 2'b10;
      13'h001a: color = 2'b11;
      13'h001b: color = 2'b11;
      13'h001c: color = 2'b11;
      13'h001d: color = 2'b11;
      13'h001e: color = 2'b11;
      13'h001f: color = 2'b11;
      13'h0020: color = 2'b11;
      13'h0021: color = 2'b11;
      13'h0022: color = 2'b00;
      13'h0023: color = 2'b00;
      13'h0024: color = 2'b00;
      13'h0025: color = 2'b00;
      13'h0026: color = 2'b00;
      13'h0027: color = 2'b00;
      13'h0028: color = 2'b00;
      13'h0029: color = 2'b00;
      13'h002a: color = 2'b00;
      13'h002b: color = 2'b00;
      13'h002c: color = 2'b00;
      13'h002d: color = 2'b00;
      13'h002e: color = 2'b00;
      13'h002f: color = 2'b00;
      13'h0030: color = 2'b00;
      13'h0031: color = 2'b00;
      13'h0032: color = 2'b00;
      13'h0033: color = 2'b00;
      13'h0034: color = 2'b00;
      13'h0035: color = 2'b00;
      13'h0036: color = 2'b00;
      13'h0037: color = 2'b00;
      13'h0038: color = 2'b00;
      13'h0039: color = 2'b00;
      13'h003a: color = 2'b00;
      13'h003b: color = 2'b00;
      13'h003c: color = 2'b00;
      13'h003d: color = 2'b00;
      13'h003e: color = 2'b00;
      13'h003f: color = 2'b00;
      13'h0040: color = 2'b00;
      13'h0041: color = 2'b00;
      13'h0042: color = 2'b00;
      13'h0043: color = 2'b00;
      13'h0044: color = 2'b00;
      13'h0045: color = 2'b00;
      13'h0046: color = 2'b00;
      13'h0047: color = 2'b00;
      13'h0048: color = 2'b00;
      13'h0049: color = 2'b00;
      13'h004a: color = 2'b00;
      13'h004b: color = 2'b00;
      13'h004c: color = 2'b00;
      13'h004d: color = 2'b00;
      13'h004e: color = 2'b00;
      13'h004f: color = 2'b00;
      13'h0050: color = 2'b00;
      13'h0051: color = 2'b00;
      13'h0052: color = 2'b00;
      13'h0053: color = 2'b00;
      13'h0054: color = 2'b00;
      13'h0055: color = 2'b00;
      13'h0056: color = 2'b00;
      13'h0057: color = 2'b00;
      13'h0058: color = 2'b00;
      13'h0059: color = 2'b00;
      13'h005a: color = 2'b00;
      13'h005b: color = 2'b00;
      13'h005c: color = 2'b00;
      13'h005d: color = 2'b00;
      13'h005e: color = 2'b11;
      13'h005f: color = 2'b11;
      13'h0060: color = 2'b11;
      13'h0061: color = 2'b11;
      13'h0062: color = 2'b11;
      13'h0063: color = 2'b11;
      13'h0064: color = 2'b10;
      13'h0065: color = 2'b10;
      13'h0066: color = 2'b11;
      13'h0067: color = 2'b11;
      13'h0068: color = 2'b10;
      13'h0069: color = 2'b10;
      13'h006a: color = 2'b11;
      13'h006b: color = 2'b11;
      13'h006c: color = 2'b11;
      13'h006d: color = 2'b11;
      13'h006e: color = 2'b11;
      13'h006f: color = 2'b11;
      13'h0070: color = 2'b11;
      13'h0071: color = 2'b11;
      13'h0072: color = 2'b11;
      13'h0073: color = 2'b11;
      13'h0074: color = 2'b10;
      13'h0075: color = 2'b10;
      13'h0076: color = 2'b11;
      13'h0077: color = 2'b11;
      13'h0078: color = 2'b10;
      13'h0079: color = 2'b10;
      13'h007a: color = 2'b11;
      13'h007b: color = 2'b11;
      13'h007c: color = 2'b11;
      13'h007d: color = 2'b11;
      13'h007e: color = 2'b11;
      13'h007f: color = 2'b11;
      13'h0080: color = 2'b11;
      13'h0081: color = 2'b11;
      13'h0082: color = 2'b11;
      13'h0083: color = 2'b11;
      13'h0084: color = 2'b10;
      13'h0085: color = 2'b10;
      13'h0086: color = 2'b11;
      13'h0087: color = 2'b11;
      13'h0088: color = 2'b10;
      13'h0089: color = 2'b10;
      13'h008a: color = 2'b11;
      13'h008b: color = 2'b11;
      13'h008c: color = 2'b11;
      13'h008d: color = 2'b11;
      13'h008e: color = 2'b11;
      13'h008f: color = 2'b11;
      13'h0090: color = 2'b11;
      13'h0091: color = 2'b11;
      13'h0092: color = 2'b11;
      13'h0093: color = 2'b11;
      13'h0094: color = 2'b10;
      13'h0095: color = 2'b10;
      13'h0096: color = 2'b11;
      13'h0097: color = 2'b11;
      13'h0098: color = 2'b10;
      13'h0099: color = 2'b10;
      13'h009a: color = 2'b11;
      13'h009b: color = 2'b11;
      13'h009c: color = 2'b11;
      13'h009d: color = 2'b11;
      13'h009e: color = 2'b11;
      13'h009f: color = 2'b11;
      13'h00a0: color = 2'b11;
      13'h00a1: color = 2'b11;
      13'h00a2: color = 2'b00;
      13'h00a3: color = 2'b00;
      13'h00a4: color = 2'b00;
      13'h00a5: color = 2'b00;
      13'h00a6: color = 2'b00;
      13'h00a7: color = 2'b00;
      13'h00a8: color = 2'b00;
      13'h00a9: color = 2'b00;
      13'h00aa: color = 2'b00;
      13'h00ab: color = 2'b00;
      13'h00ac: color = 2'b00;
      13'h00ad: color = 2'b00;
      13'h00ae: color = 2'b00;
      13'h00af: color = 2'b00;
      13'h00b0: color = 2'b00;
      13'h00b1: color = 2'b00;
      13'h00b2: color = 2'b00;
      13'h00b3: color = 2'b00;
      13'h00b4: color = 2'b00;
      13'h00b5: color = 2'b00;
      13'h00b6: color = 2'b00;
      13'h00b7: color = 2'b00;
      13'h00b8: color = 2'b00;
      13'h00b9: color = 2'b00;
      13'h00ba: color = 2'b00;
      13'h00bb: color = 2'b00;
      13'h00bc: color = 2'b00;
      13'h00bd: color = 2'b00;
      13'h00be: color = 2'b00;
      13'h00bf: color = 2'b00;
      13'h00c0: color = 2'b00;
      13'h00c1: color = 2'b00;
      13'h00c2: color = 2'b00;
      13'h00c3: color = 2'b00;
      13'h00c4: color = 2'b00;
      13'h00c5: color = 2'b00;
      13'h00c6: color = 2'b00;
      13'h00c7: color = 2'b00;
      13'h00c8: color = 2'b00;
      13'h00c9: color = 2'b00;
      13'h00ca: color = 2'b00;
      13'h00cb: color = 2'b00;
      13'h00cc: color = 2'b00;
      13'h00cd: color = 2'b00;
      13'h00ce: color = 2'b00;
      13'h00cf: color = 2'b00;
      13'h00d0: color = 2'b00;
      13'h00d1: color = 2'b00;
      13'h00d2: color = 2'b00;
      13'h00d3: color = 2'b00;
      13'h00d4: color = 2'b00;
      13'h00d5: color = 2'b00;
      13'h00d6: color = 2'b00;
      13'h00d7: color = 2'b00;
      13'h00d8: color = 2'b00;
      13'h00d9: color = 2'b00;
      13'h00da: color = 2'b00;
      13'h00db: color = 2'b00;
      13'h00dc: color = 2'b00;
      13'h00dd: color = 2'b00;
      13'h00de: color = 2'b11;
      13'h00df: color = 2'b11;
      13'h00e0: color = 2'b11;
      13'h00e1: color = 2'b11;
      13'h00e2: color = 2'b11;
      13'h00e3: color = 2'b11;
      13'h00e4: color = 2'b10;
      13'h00e5: color = 2'b10;
      13'h00e6: color = 2'b11;
      13'h00e7: color = 2'b11;
      13'h00e8: color = 2'b10;
      13'h00e9: color = 2'b10;
      13'h00ea: color = 2'b11;
      13'h00eb: color = 2'b11;
      13'h00ec: color = 2'b11;
      13'h00ed: color = 2'b11;
      13'h00ee: color = 2'b11;
      13'h00ef: color = 2'b11;
      13'h00f0: color = 2'b11;
      13'h00f1: color = 2'b11;
      13'h00f2: color = 2'b11;
      13'h00f3: color = 2'b11;
      13'h00f4: color = 2'b10;
      13'h00f5: color = 2'b10;
      13'h00f6: color = 2'b11;
      13'h00f7: color = 2'b11;
      13'h00f8: color = 2'b10;
      13'h00f9: color = 2'b10;
      13'h00fa: color = 2'b11;
      13'h00fb: color = 2'b11;
      13'h00fc: color = 2'b11;
      13'h00fd: color = 2'b11;
      13'h00fe: color = 2'b11;
      13'h00ff: color = 2'b11;
      13'h0100: color = 2'b11;
      13'h0101: color = 2'b11;
      13'h0102: color = 2'b10;
      13'h0103: color = 2'b10;
      13'h0104: color = 2'b11;
      13'h0105: color = 2'b11;
      13'h0106: color = 2'b11;
      13'h0107: color = 2'b11;
      13'h0108: color = 2'b11;
      13'h0109: color = 2'b11;
      13'h010a: color = 2'b10;
      13'h010b: color = 2'b10;
      13'h010c: color = 2'b11;
      13'h010d: color = 2'b11;
      13'h010e: color = 2'b11;
      13'h010f: color = 2'b11;
      13'h0110: color = 2'b11;
      13'h0111: color = 2'b11;
      13'h0112: color = 2'b10;
      13'h0113: color = 2'b10;
      13'h0114: color = 2'b11;
      13'h0115: color = 2'b11;
      13'h0116: color = 2'b11;
      13'h0117: color = 2'b11;
      13'h0118: color = 2'b11;
      13'h0119: color = 2'b11;
      13'h011a: color = 2'b10;
      13'h011b: color = 2'b10;
      13'h011c: color = 2'b11;
      13'h011d: color = 2'b11;
      13'h011e: color = 2'b11;
      13'h011f: color = 2'b11;
      13'h0120: color = 2'b00;
      13'h0121: color = 2'b00;
      13'h0122: color = 2'b11;
      13'h0123: color = 2'b11;
      13'h0124: color = 2'b11;
      13'h0125: color = 2'b11;
      13'h0126: color = 2'b11;
      13'h0127: color = 2'b11;
      13'h0128: color = 2'b11;
      13'h0129: color = 2'b11;
      13'h012a: color = 2'b11;
      13'h012b: color = 2'b11;
      13'h012c: color = 2'b11;
      13'h012d: color = 2'b11;
      13'h012e: color = 2'b11;
      13'h012f: color = 2'b11;
      13'h0130: color = 2'b11;
      13'h0131: color = 2'b11;
      13'h0132: color = 2'b11;
      13'h0133: color = 2'b11;
      13'h0134: color = 2'b11;
      13'h0135: color = 2'b11;
      13'h0136: color = 2'b11;
      13'h0137: color = 2'b11;
      13'h0138: color = 2'b11;
      13'h0139: color = 2'b11;
      13'h013a: color = 2'b11;
      13'h013b: color = 2'b11;
      13'h013c: color = 2'b11;
      13'h013d: color = 2'b11;
      13'h013e: color = 2'b11;
      13'h013f: color = 2'b11;
      13'h0140: color = 2'b11;
      13'h0141: color = 2'b11;
      13'h0142: color = 2'b11;
      13'h0143: color = 2'b11;
      13'h0144: color = 2'b11;
      13'h0145: color = 2'b11;
      13'h0146: color = 2'b11;
      13'h0147: color = 2'b11;
      13'h0148: color = 2'b11;
      13'h0149: color = 2'b11;
      13'h014a: color = 2'b11;
      13'h014b: color = 2'b11;
      13'h014c: color = 2'b11;
      13'h014d: color = 2'b11;
      13'h014e: color = 2'b11;
      13'h014f: color = 2'b11;
      13'h0150: color = 2'b11;
      13'h0151: color = 2'b11;
      13'h0152: color = 2'b11;
      13'h0153: color = 2'b11;
      13'h0154: color = 2'b11;
      13'h0155: color = 2'b11;
      13'h0156: color = 2'b11;
      13'h0157: color = 2'b11;
      13'h0158: color = 2'b11;
      13'h0159: color = 2'b11;
      13'h015a: color = 2'b11;
      13'h015b: color = 2'b11;
      13'h015c: color = 2'b11;
      13'h015d: color = 2'b11;
      13'h015e: color = 2'b00;
      13'h015f: color = 2'b00;
      13'h0160: color = 2'b11;
      13'h0161: color = 2'b11;
      13'h0162: color = 2'b10;
      13'h0163: color = 2'b10;
      13'h0164: color = 2'b11;
      13'h0165: color = 2'b11;
      13'h0166: color = 2'b11;
      13'h0167: color = 2'b11;
      13'h0168: color = 2'b11;
      13'h0169: color = 2'b11;
      13'h016a: color = 2'b10;
      13'h016b: color = 2'b10;
      13'h016c: color = 2'b11;
      13'h016d: color = 2'b11;
      13'h016e: color = 2'b11;
      13'h016f: color = 2'b11;
      13'h0170: color = 2'b11;
      13'h0171: color = 2'b11;
      13'h0172: color = 2'b10;
      13'h0173: color = 2'b10;
      13'h0174: color = 2'b11;
      13'h0175: color = 2'b11;
      13'h0176: color = 2'b11;
      13'h0177: color = 2'b11;
      13'h0178: color = 2'b11;
      13'h0179: color = 2'b11;
      13'h017a: color = 2'b10;
      13'h017b: color = 2'b10;
      13'h017c: color = 2'b11;
      13'h017d: color = 2'b11;
      13'h017e: color = 2'b11;
      13'h017f: color = 2'b11;
      13'h0180: color = 2'b11;
      13'h0181: color = 2'b11;
      13'h0182: color = 2'b10;
      13'h0183: color = 2'b10;
      13'h0184: color = 2'b11;
      13'h0185: color = 2'b11;
      13'h0186: color = 2'b11;
      13'h0187: color = 2'b11;
      13'h0188: color = 2'b11;
      13'h0189: color = 2'b11;
      13'h018a: color = 2'b10;
      13'h018b: color = 2'b10;
      13'h018c: color = 2'b11;
      13'h018d: color = 2'b11;
      13'h018e: color = 2'b11;
      13'h018f: color = 2'b11;
      13'h0190: color = 2'b11;
      13'h0191: color = 2'b11;
      13'h0192: color = 2'b10;
      13'h0193: color = 2'b10;
      13'h0194: color = 2'b11;
      13'h0195: color = 2'b11;
      13'h0196: color = 2'b11;
      13'h0197: color = 2'b11;
      13'h0198: color = 2'b11;
      13'h0199: color = 2'b11;
      13'h019a: color = 2'b10;
      13'h019b: color = 2'b10;
      13'h019c: color = 2'b11;
      13'h019d: color = 2'b11;
      13'h019e: color = 2'b11;
      13'h019f: color = 2'b11;
      13'h01a0: color = 2'b00;
      13'h01a1: color = 2'b00;
      13'h01a2: color = 2'b11;
      13'h01a3: color = 2'b11;
      13'h01a4: color = 2'b11;
      13'h01a5: color = 2'b11;
      13'h01a6: color = 2'b11;
      13'h01a7: color = 2'b11;
      13'h01a8: color = 2'b11;
      13'h01a9: color = 2'b11;
      13'h01aa: color = 2'b11;
      13'h01ab: color = 2'b11;
      13'h01ac: color = 2'b11;
      13'h01ad: color = 2'b11;
      13'h01ae: color = 2'b11;
      13'h01af: color = 2'b11;
      13'h01b0: color = 2'b11;
      13'h01b1: color = 2'b11;
      13'h01b2: color = 2'b11;
      13'h01b3: color = 2'b11;
      13'h01b4: color = 2'b11;
      13'h01b5: color = 2'b11;
      13'h01b6: color = 2'b11;
      13'h01b7: color = 2'b11;
      13'h01b8: color = 2'b11;
      13'h01b9: color = 2'b11;
      13'h01ba: color = 2'b11;
      13'h01bb: color = 2'b11;
      13'h01bc: color = 2'b11;
      13'h01bd: color = 2'b11;
      13'h01be: color = 2'b11;
      13'h01bf: color = 2'b11;
      13'h01c0: color = 2'b11;
      13'h01c1: color = 2'b11;
      13'h01c2: color = 2'b11;
      13'h01c3: color = 2'b11;
      13'h01c4: color = 2'b11;
      13'h01c5: color = 2'b11;
      13'h01c6: color = 2'b11;
      13'h01c7: color = 2'b11;
      13'h01c8: color = 2'b11;
      13'h01c9: color = 2'b11;
      13'h01ca: color = 2'b11;
      13'h01cb: color = 2'b11;
      13'h01cc: color = 2'b11;
      13'h01cd: color = 2'b11;
      13'h01ce: color = 2'b11;
      13'h01cf: color = 2'b11;
      13'h01d0: color = 2'b11;
      13'h01d1: color = 2'b11;
      13'h01d2: color = 2'b11;
      13'h01d3: color = 2'b11;
      13'h01d4: color = 2'b11;
      13'h01d5: color = 2'b11;
      13'h01d6: color = 2'b11;
      13'h01d7: color = 2'b11;
      13'h01d8: color = 2'b11;
      13'h01d9: color = 2'b11;
      13'h01da: color = 2'b11;
      13'h01db: color = 2'b11;
      13'h01dc: color = 2'b11;
      13'h01dd: color = 2'b11;
      13'h01de: color = 2'b00;
      13'h01df: color = 2'b00;
      13'h01e0: color = 2'b11;
      13'h01e1: color = 2'b11;
      13'h01e2: color = 2'b10;
      13'h01e3: color = 2'b10;
      13'h01e4: color = 2'b11;
      13'h01e5: color = 2'b11;
      13'h01e6: color = 2'b11;
      13'h01e7: color = 2'b11;
      13'h01e8: color = 2'b11;
      13'h01e9: color = 2'b11;
      13'h01ea: color = 2'b10;
      13'h01eb: color = 2'b10;
      13'h01ec: color = 2'b11;
      13'h01ed: color = 2'b11;
      13'h01ee: color = 2'b11;
      13'h01ef: color = 2'b11;
      13'h01f0: color = 2'b11;
      13'h01f1: color = 2'b11;
      13'h01f2: color = 2'b10;
      13'h01f3: color = 2'b10;
      13'h01f4: color = 2'b11;
      13'h01f5: color = 2'b11;
      13'h01f6: color = 2'b11;
      13'h01f7: color = 2'b11;
      13'h01f8: color = 2'b11;
      13'h01f9: color = 2'b11;
      13'h01fa: color = 2'b10;
      13'h01fb: color = 2'b10;
      13'h01fc: color = 2'b11;
      13'h01fd: color = 2'b11;
      13'h01fe: color = 2'b11;
      13'h01ff: color = 2'b11;
      13'h0200: color = 2'b10;
      13'h0201: color = 2'b10;
      13'h0202: color = 2'b11;
      13'h0203: color = 2'b11;
      13'h0204: color = 2'b11;
      13'h0205: color = 2'b11;
      13'h0206: color = 2'b11;
      13'h0207: color = 2'b11;
      13'h0208: color = 2'b11;
      13'h0209: color = 2'b11;
      13'h020a: color = 2'b11;
      13'h020b: color = 2'b11;
      13'h020c: color = 2'b10;
      13'h020d: color = 2'b10;
      13'h020e: color = 2'b11;
      13'h020f: color = 2'b11;
      13'h0210: color = 2'b10;
      13'h0211: color = 2'b10;
      13'h0212: color = 2'b11;
      13'h0213: color = 2'b11;
      13'h0214: color = 2'b11;
      13'h0215: color = 2'b11;
      13'h0216: color = 2'b11;
      13'h0217: color = 2'b11;
      13'h0218: color = 2'b11;
      13'h0219: color = 2'b11;
      13'h021a: color = 2'b11;
      13'h021b: color = 2'b11;
      13'h021c: color = 2'b10;
      13'h021d: color = 2'b10;
      13'h021e: color = 2'b11;
      13'h021f: color = 2'b11;
      13'h0220: color = 2'b00;
      13'h0221: color = 2'b00;
      13'h0222: color = 2'b11;
      13'h0223: color = 2'b11;
      13'h0224: color = 2'b10;
      13'h0225: color = 2'b10;
      13'h0226: color = 2'b10;
      13'h0227: color = 2'b10;
      13'h0228: color = 2'b10;
      13'h0229: color = 2'b10;
      13'h022a: color = 2'b10;
      13'h022b: color = 2'b10;
      13'h022c: color = 2'b10;
      13'h022d: color = 2'b10;
      13'h022e: color = 2'b10;
      13'h022f: color = 2'b10;
      13'h0230: color = 2'b10;
      13'h0231: color = 2'b10;
      13'h0232: color = 2'b10;
      13'h0233: color = 2'b10;
      13'h0234: color = 2'b10;
      13'h0235: color = 2'b10;
      13'h0236: color = 2'b10;
      13'h0237: color = 2'b10;
      13'h0238: color = 2'b10;
      13'h0239: color = 2'b10;
      13'h023a: color = 2'b10;
      13'h023b: color = 2'b10;
      13'h023c: color = 2'b10;
      13'h023d: color = 2'b10;
      13'h023e: color = 2'b10;
      13'h023f: color = 2'b10;
      13'h0240: color = 2'b10;
      13'h0241: color = 2'b10;
      13'h0242: color = 2'b10;
      13'h0243: color = 2'b10;
      13'h0244: color = 2'b10;
      13'h0245: color = 2'b10;
      13'h0246: color = 2'b10;
      13'h0247: color = 2'b10;
      13'h0248: color = 2'b10;
      13'h0249: color = 2'b10;
      13'h024a: color = 2'b10;
      13'h024b: color = 2'b10;
      13'h024c: color = 2'b10;
      13'h024d: color = 2'b10;
      13'h024e: color = 2'b10;
      13'h024f: color = 2'b10;
      13'h0250: color = 2'b10;
      13'h0251: color = 2'b10;
      13'h0252: color = 2'b10;
      13'h0253: color = 2'b10;
      13'h0254: color = 2'b10;
      13'h0255: color = 2'b10;
      13'h0256: color = 2'b10;
      13'h0257: color = 2'b10;
      13'h0258: color = 2'b10;
      13'h0259: color = 2'b10;
      13'h025a: color = 2'b10;
      13'h025b: color = 2'b10;
      13'h025c: color = 2'b01;
      13'h025d: color = 2'b01;
      13'h025e: color = 2'b00;
      13'h025f: color = 2'b00;
      13'h0260: color = 2'b10;
      13'h0261: color = 2'b10;
      13'h0262: color = 2'b11;
      13'h0263: color = 2'b11;
      13'h0264: color = 2'b11;
      13'h0265: color = 2'b11;
      13'h0266: color = 2'b11;
      13'h0267: color = 2'b11;
      13'h0268: color = 2'b11;
      13'h0269: color = 2'b11;
      13'h026a: color = 2'b11;
      13'h026b: color = 2'b11;
      13'h026c: color = 2'b10;
      13'h026d: color = 2'b10;
      13'h026e: color = 2'b11;
      13'h026f: color = 2'b11;
      13'h0270: color = 2'b10;
      13'h0271: color = 2'b10;
      13'h0272: color = 2'b11;
      13'h0273: color = 2'b11;
      13'h0274: color = 2'b11;
      13'h0275: color = 2'b11;
      13'h0276: color = 2'b11;
      13'h0277: color = 2'b11;
      13'h0278: color = 2'b11;
      13'h0279: color = 2'b11;
      13'h027a: color = 2'b11;
      13'h027b: color = 2'b11;
      13'h027c: color = 2'b10;
      13'h027d: color = 2'b10;
      13'h027e: color = 2'b11;
      13'h027f: color = 2'b11;
      13'h0280: color = 2'b10;
      13'h0281: color = 2'b10;
      13'h0282: color = 2'b11;
      13'h0283: color = 2'b11;
      13'h0284: color = 2'b11;
      13'h0285: color = 2'b11;
      13'h0286: color = 2'b11;
      13'h0287: color = 2'b11;
      13'h0288: color = 2'b11;
      13'h0289: color = 2'b11;
      13'h028a: color = 2'b11;
      13'h028b: color = 2'b11;
      13'h028c: color = 2'b10;
      13'h028d: color = 2'b10;
      13'h028e: color = 2'b11;
      13'h028f: color = 2'b11;
      13'h0290: color = 2'b10;
      13'h0291: color = 2'b10;
      13'h0292: color = 2'b11;
      13'h0293: color = 2'b11;
      13'h0294: color = 2'b11;
      13'h0295: color = 2'b11;
      13'h0296: color = 2'b11;
      13'h0297: color = 2'b11;
      13'h0298: color = 2'b11;
      13'h0299: color = 2'b11;
      13'h029a: color = 2'b11;
      13'h029b: color = 2'b11;
      13'h029c: color = 2'b10;
      13'h029d: color = 2'b10;
      13'h029e: color = 2'b11;
      13'h029f: color = 2'b11;
      13'h02a0: color = 2'b00;
      13'h02a1: color = 2'b00;
      13'h02a2: color = 2'b11;
      13'h02a3: color = 2'b11;
      13'h02a4: color = 2'b10;
      13'h02a5: color = 2'b10;
      13'h02a6: color = 2'b10;
      13'h02a7: color = 2'b10;
      13'h02a8: color = 2'b10;
      13'h02a9: color = 2'b10;
      13'h02aa: color = 2'b10;
      13'h02ab: color = 2'b10;
      13'h02ac: color = 2'b10;
      13'h02ad: color = 2'b10;
      13'h02ae: color = 2'b10;
      13'h02af: color = 2'b10;
      13'h02b0: color = 2'b10;
      13'h02b1: color = 2'b10;
      13'h02b2: color = 2'b10;
      13'h02b3: color = 2'b10;
      13'h02b4: color = 2'b10;
      13'h02b5: color = 2'b10;
      13'h02b6: color = 2'b10;
      13'h02b7: color = 2'b10;
      13'h02b8: color = 2'b10;
      13'h02b9: color = 2'b10;
      13'h02ba: color = 2'b10;
      13'h02bb: color = 2'b10;
      13'h02bc: color = 2'b10;
      13'h02bd: color = 2'b10;
      13'h02be: color = 2'b10;
      13'h02bf: color = 2'b10;
      13'h02c0: color = 2'b10;
      13'h02c1: color = 2'b10;
      13'h02c2: color = 2'b10;
      13'h02c3: color = 2'b10;
      13'h02c4: color = 2'b10;
      13'h02c5: color = 2'b10;
      13'h02c6: color = 2'b10;
      13'h02c7: color = 2'b10;
      13'h02c8: color = 2'b10;
      13'h02c9: color = 2'b10;
      13'h02ca: color = 2'b10;
      13'h02cb: color = 2'b10;
      13'h02cc: color = 2'b10;
      13'h02cd: color = 2'b10;
      13'h02ce: color = 2'b10;
      13'h02cf: color = 2'b10;
      13'h02d0: color = 2'b10;
      13'h02d1: color = 2'b10;
      13'h02d2: color = 2'b10;
      13'h02d3: color = 2'b10;
      13'h02d4: color = 2'b10;
      13'h02d5: color = 2'b10;
      13'h02d6: color = 2'b10;
      13'h02d7: color = 2'b10;
      13'h02d8: color = 2'b10;
      13'h02d9: color = 2'b10;
      13'h02da: color = 2'b10;
      13'h02db: color = 2'b10;
      13'h02dc: color = 2'b01;
      13'h02dd: color = 2'b01;
      13'h02de: color = 2'b00;
      13'h02df: color = 2'b00;
      13'h02e0: color = 2'b10;
      13'h02e1: color = 2'b10;
      13'h02e2: color = 2'b11;
      13'h02e3: color = 2'b11;
      13'h02e4: color = 2'b11;
      13'h02e5: color = 2'b11;
      13'h02e6: color = 2'b11;
      13'h02e7: color = 2'b11;
      13'h02e8: color = 2'b11;
      13'h02e9: color = 2'b11;
      13'h02ea: color = 2'b11;
      13'h02eb: color = 2'b11;
      13'h02ec: color = 2'b10;
      13'h02ed: color = 2'b10;
      13'h02ee: color = 2'b11;
      13'h02ef: color = 2'b11;
      13'h02f0: color = 2'b10;
      13'h02f1: color = 2'b10;
      13'h02f2: color = 2'b11;
      13'h02f3: color = 2'b11;
      13'h02f4: color = 2'b11;
      13'h02f5: color = 2'b11;
      13'h02f6: color = 2'b11;
      13'h02f7: color = 2'b11;
      13'h02f8: color = 2'b11;
      13'h02f9: color = 2'b11;
      13'h02fa: color = 2'b11;
      13'h02fb: color = 2'b11;
      13'h02fc: color = 2'b10;
      13'h02fd: color = 2'b10;
      13'h02fe: color = 2'b11;
      13'h02ff: color = 2'b11;
      13'h0300: color = 2'b11;
      13'h0301: color = 2'b11;
      13'h0302: color = 2'b11;
      13'h0303: color = 2'b11;
      13'h0304: color = 2'b11;
      13'h0305: color = 2'b11;
      13'h0306: color = 2'b11;
      13'h0307: color = 2'b11;
      13'h0308: color = 2'b11;
      13'h0309: color = 2'b11;
      13'h030a: color = 2'b11;
      13'h030b: color = 2'b11;
      13'h030c: color = 2'b11;
      13'h030d: color = 2'b11;
      13'h030e: color = 2'b10;
      13'h030f: color = 2'b10;
      13'h0310: color = 2'b11;
      13'h0311: color = 2'b11;
      13'h0312: color = 2'b11;
      13'h0313: color = 2'b11;
      13'h0314: color = 2'b11;
      13'h0315: color = 2'b11;
      13'h0316: color = 2'b11;
      13'h0317: color = 2'b11;
      13'h0318: color = 2'b11;
      13'h0319: color = 2'b11;
      13'h031a: color = 2'b11;
      13'h031b: color = 2'b11;
      13'h031c: color = 2'b11;
      13'h031d: color = 2'b11;
      13'h031e: color = 2'b10;
      13'h031f: color = 2'b10;
      13'h0320: color = 2'b00;
      13'h0321: color = 2'b00;
      13'h0322: color = 2'b11;
      13'h0323: color = 2'b11;
      13'h0324: color = 2'b10;
      13'h0325: color = 2'b10;
      13'h0326: color = 2'b10;
      13'h0327: color = 2'b10;
      13'h0328: color = 2'b10;
      13'h0329: color = 2'b10;
      13'h032a: color = 2'b10;
      13'h032b: color = 2'b10;
      13'h032c: color = 2'b10;
      13'h032d: color = 2'b10;
      13'h032e: color = 2'b10;
      13'h032f: color = 2'b10;
      13'h0330: color = 2'b10;
      13'h0331: color = 2'b10;
      13'h0332: color = 2'b10;
      13'h0333: color = 2'b10;
      13'h0334: color = 2'b10;
      13'h0335: color = 2'b10;
      13'h0336: color = 2'b10;
      13'h0337: color = 2'b10;
      13'h0338: color = 2'b10;
      13'h0339: color = 2'b10;
      13'h033a: color = 2'b10;
      13'h033b: color = 2'b10;
      13'h033c: color = 2'b10;
      13'h033d: color = 2'b10;
      13'h033e: color = 2'b10;
      13'h033f: color = 2'b10;
      13'h0340: color = 2'b10;
      13'h0341: color = 2'b10;
      13'h0342: color = 2'b10;
      13'h0343: color = 2'b10;
      13'h0344: color = 2'b10;
      13'h0345: color = 2'b10;
      13'h0346: color = 2'b10;
      13'h0347: color = 2'b10;
      13'h0348: color = 2'b10;
      13'h0349: color = 2'b10;
      13'h034a: color = 2'b10;
      13'h034b: color = 2'b10;
      13'h034c: color = 2'b10;
      13'h034d: color = 2'b10;
      13'h034e: color = 2'b10;
      13'h034f: color = 2'b10;
      13'h0350: color = 2'b10;
      13'h0351: color = 2'b10;
      13'h0352: color = 2'b10;
      13'h0353: color = 2'b10;
      13'h0354: color = 2'b10;
      13'h0355: color = 2'b10;
      13'h0356: color = 2'b10;
      13'h0357: color = 2'b10;
      13'h0358: color = 2'b10;
      13'h0359: color = 2'b10;
      13'h035a: color = 2'b10;
      13'h035b: color = 2'b10;
      13'h035c: color = 2'b01;
      13'h035d: color = 2'b01;
      13'h035e: color = 2'b00;
      13'h035f: color = 2'b00;
      13'h0360: color = 2'b11;
      13'h0361: color = 2'b11;
      13'h0362: color = 2'b11;
      13'h0363: color = 2'b11;
      13'h0364: color = 2'b11;
      13'h0365: color = 2'b11;
      13'h0366: color = 2'b11;
      13'h0367: color = 2'b11;
      13'h0368: color = 2'b11;
      13'h0369: color = 2'b11;
      13'h036a: color = 2'b11;
      13'h036b: color = 2'b11;
      13'h036c: color = 2'b11;
      13'h036d: color = 2'b11;
      13'h036e: color = 2'b10;
      13'h036f: color = 2'b10;
      13'h0370: color = 2'b11;
      13'h0371: color = 2'b11;
      13'h0372: color = 2'b11;
      13'h0373: color = 2'b11;
      13'h0374: color = 2'b11;
      13'h0375: color = 2'b11;
      13'h0376: color = 2'b11;
      13'h0377: color = 2'b11;
      13'h0378: color = 2'b11;
      13'h0379: color = 2'b11;
      13'h037a: color = 2'b11;
      13'h037b: color = 2'b11;
      13'h037c: color = 2'b11;
      13'h037d: color = 2'b11;
      13'h037e: color = 2'b10;
      13'h037f: color = 2'b10;
      13'h0380: color = 2'b11;
      13'h0381: color = 2'b11;
      13'h0382: color = 2'b11;
      13'h0383: color = 2'b11;
      13'h0384: color = 2'b11;
      13'h0385: color = 2'b11;
      13'h0386: color = 2'b11;
      13'h0387: color = 2'b11;
      13'h0388: color = 2'b11;
      13'h0389: color = 2'b11;
      13'h038a: color = 2'b11;
      13'h038b: color = 2'b11;
      13'h038c: color = 2'b11;
      13'h038d: color = 2'b11;
      13'h038e: color = 2'b10;
      13'h038f: color = 2'b10;
      13'h0390: color = 2'b11;
      13'h0391: color = 2'b11;
      13'h0392: color = 2'b11;
      13'h0393: color = 2'b11;
      13'h0394: color = 2'b11;
      13'h0395: color = 2'b11;
      13'h0396: color = 2'b11;
      13'h0397: color = 2'b11;
      13'h0398: color = 2'b11;
      13'h0399: color = 2'b11;
      13'h039a: color = 2'b11;
      13'h039b: color = 2'b11;
      13'h039c: color = 2'b11;
      13'h039d: color = 2'b11;
      13'h039e: color = 2'b10;
      13'h039f: color = 2'b10;
      13'h03a0: color = 2'b00;
      13'h03a1: color = 2'b00;
      13'h03a2: color = 2'b11;
      13'h03a3: color = 2'b11;
      13'h03a4: color = 2'b10;
      13'h03a5: color = 2'b10;
      13'h03a6: color = 2'b10;
      13'h03a7: color = 2'b10;
      13'h03a8: color = 2'b10;
      13'h03a9: color = 2'b10;
      13'h03aa: color = 2'b10;
      13'h03ab: color = 2'b10;
      13'h03ac: color = 2'b10;
      13'h03ad: color = 2'b10;
      13'h03ae: color = 2'b10;
      13'h03af: color = 2'b10;
      13'h03b0: color = 2'b10;
      13'h03b1: color = 2'b10;
      13'h03b2: color = 2'b10;
      13'h03b3: color = 2'b10;
      13'h03b4: color = 2'b10;
      13'h03b5: color = 2'b10;
      13'h03b6: color = 2'b10;
      13'h03b7: color = 2'b10;
      13'h03b8: color = 2'b10;
      13'h03b9: color = 2'b10;
      13'h03ba: color = 2'b10;
      13'h03bb: color = 2'b10;
      13'h03bc: color = 2'b10;
      13'h03bd: color = 2'b10;
      13'h03be: color = 2'b10;
      13'h03bf: color = 2'b10;
      13'h03c0: color = 2'b10;
      13'h03c1: color = 2'b10;
      13'h03c2: color = 2'b10;
      13'h03c3: color = 2'b10;
      13'h03c4: color = 2'b10;
      13'h03c5: color = 2'b10;
      13'h03c6: color = 2'b10;
      13'h03c7: color = 2'b10;
      13'h03c8: color = 2'b10;
      13'h03c9: color = 2'b10;
      13'h03ca: color = 2'b10;
      13'h03cb: color = 2'b10;
      13'h03cc: color = 2'b10;
      13'h03cd: color = 2'b10;
      13'h03ce: color = 2'b10;
      13'h03cf: color = 2'b10;
      13'h03d0: color = 2'b10;
      13'h03d1: color = 2'b10;
      13'h03d2: color = 2'b10;
      13'h03d3: color = 2'b10;
      13'h03d4: color = 2'b10;
      13'h03d5: color = 2'b10;
      13'h03d6: color = 2'b10;
      13'h03d7: color = 2'b10;
      13'h03d8: color = 2'b10;
      13'h03d9: color = 2'b10;
      13'h03da: color = 2'b10;
      13'h03db: color = 2'b10;
      13'h03dc: color = 2'b01;
      13'h03dd: color = 2'b01;
      13'h03de: color = 2'b00;
      13'h03df: color = 2'b00;
      13'h03e0: color = 2'b11;
      13'h03e1: color = 2'b11;
      13'h03e2: color = 2'b11;
      13'h03e3: color = 2'b11;
      13'h03e4: color = 2'b11;
      13'h03e5: color = 2'b11;
      13'h03e6: color = 2'b11;
      13'h03e7: color = 2'b11;
      13'h03e8: color = 2'b11;
      13'h03e9: color = 2'b11;
      13'h03ea: color = 2'b11;
      13'h03eb: color = 2'b11;
      13'h03ec: color = 2'b11;
      13'h03ed: color = 2'b11;
      13'h03ee: color = 2'b10;
      13'h03ef: color = 2'b10;
      13'h03f0: color = 2'b11;
      13'h03f1: color = 2'b11;
      13'h03f2: color = 2'b11;
      13'h03f3: color = 2'b11;
      13'h03f4: color = 2'b11;
      13'h03f5: color = 2'b11;
      13'h03f6: color = 2'b11;
      13'h03f7: color = 2'b11;
      13'h03f8: color = 2'b11;
      13'h03f9: color = 2'b11;
      13'h03fa: color = 2'b11;
      13'h03fb: color = 2'b11;
      13'h03fc: color = 2'b11;
      13'h03fd: color = 2'b11;
      13'h03fe: color = 2'b10;
      13'h03ff: color = 2'b10;
      13'h0400: color = 2'b10;
      13'h0401: color = 2'b10;
      13'h0402: color = 2'b11;
      13'h0403: color = 2'b11;
      13'h0404: color = 2'b11;
      13'h0405: color = 2'b11;
      13'h0406: color = 2'b11;
      13'h0407: color = 2'b11;
      13'h0408: color = 2'b11;
      13'h0409: color = 2'b11;
      13'h040a: color = 2'b11;
      13'h040b: color = 2'b11;
      13'h040c: color = 2'b11;
      13'h040d: color = 2'b11;
      13'h040e: color = 2'b11;
      13'h040f: color = 2'b11;
      13'h0410: color = 2'b10;
      13'h0411: color = 2'b10;
      13'h0412: color = 2'b11;
      13'h0413: color = 2'b11;
      13'h0414: color = 2'b11;
      13'h0415: color = 2'b11;
      13'h0416: color = 2'b11;
      13'h0417: color = 2'b11;
      13'h0418: color = 2'b11;
      13'h0419: color = 2'b11;
      13'h041a: color = 2'b11;
      13'h041b: color = 2'b11;
      13'h041c: color = 2'b11;
      13'h041d: color = 2'b11;
      13'h041e: color = 2'b11;
      13'h041f: color = 2'b11;
      13'h0420: color = 2'b00;
      13'h0421: color = 2'b00;
      13'h0422: color = 2'b11;
      13'h0423: color = 2'b11;
      13'h0424: color = 2'b10;
      13'h0425: color = 2'b10;
      13'h0426: color = 2'b10;
      13'h0427: color = 2'b10;
      13'h0428: color = 2'b10;
      13'h0429: color = 2'b10;
      13'h042a: color = 2'b10;
      13'h042b: color = 2'b10;
      13'h042c: color = 2'b10;
      13'h042d: color = 2'b10;
      13'h042e: color = 2'b10;
      13'h042f: color = 2'b10;
      13'h0430: color = 2'b10;
      13'h0431: color = 2'b10;
      13'h0432: color = 2'b10;
      13'h0433: color = 2'b10;
      13'h0434: color = 2'b10;
      13'h0435: color = 2'b10;
      13'h0436: color = 2'b10;
      13'h0437: color = 2'b10;
      13'h0438: color = 2'b10;
      13'h0439: color = 2'b10;
      13'h043a: color = 2'b10;
      13'h043b: color = 2'b10;
      13'h043c: color = 2'b10;
      13'h043d: color = 2'b10;
      13'h043e: color = 2'b10;
      13'h043f: color = 2'b10;
      13'h0440: color = 2'b10;
      13'h0441: color = 2'b10;
      13'h0442: color = 2'b10;
      13'h0443: color = 2'b10;
      13'h0444: color = 2'b10;
      13'h0445: color = 2'b10;
      13'h0446: color = 2'b10;
      13'h0447: color = 2'b10;
      13'h0448: color = 2'b10;
      13'h0449: color = 2'b10;
      13'h044a: color = 2'b10;
      13'h044b: color = 2'b10;
      13'h044c: color = 2'b10;
      13'h044d: color = 2'b10;
      13'h044e: color = 2'b10;
      13'h044f: color = 2'b10;
      13'h0450: color = 2'b10;
      13'h0451: color = 2'b10;
      13'h0452: color = 2'b10;
      13'h0453: color = 2'b10;
      13'h0454: color = 2'b10;
      13'h0455: color = 2'b10;
      13'h0456: color = 2'b10;
      13'h0457: color = 2'b10;
      13'h0458: color = 2'b10;
      13'h0459: color = 2'b10;
      13'h045a: color = 2'b10;
      13'h045b: color = 2'b10;
      13'h045c: color = 2'b01;
      13'h045d: color = 2'b01;
      13'h045e: color = 2'b00;
      13'h045f: color = 2'b00;
      13'h0460: color = 2'b10;
      13'h0461: color = 2'b10;
      13'h0462: color = 2'b11;
      13'h0463: color = 2'b11;
      13'h0464: color = 2'b11;
      13'h0465: color = 2'b11;
      13'h0466: color = 2'b11;
      13'h0467: color = 2'b11;
      13'h0468: color = 2'b11;
      13'h0469: color = 2'b11;
      13'h046a: color = 2'b11;
      13'h046b: color = 2'b11;
      13'h046c: color = 2'b11;
      13'h046d: color = 2'b11;
      13'h046e: color = 2'b11;
      13'h046f: color = 2'b11;
      13'h0470: color = 2'b10;
      13'h0471: color = 2'b10;
      13'h0472: color = 2'b11;
      13'h0473: color = 2'b11;
      13'h0474: color = 2'b11;
      13'h0475: color = 2'b11;
      13'h0476: color = 2'b11;
      13'h0477: color = 2'b11;
      13'h0478: color = 2'b11;
      13'h0479: color = 2'b11;
      13'h047a: color = 2'b11;
      13'h047b: color = 2'b11;
      13'h047c: color = 2'b11;
      13'h047d: color = 2'b11;
      13'h047e: color = 2'b11;
      13'h047f: color = 2'b11;
      13'h0480: color = 2'b10;
      13'h0481: color = 2'b10;
      13'h0482: color = 2'b11;
      13'h0483: color = 2'b11;
      13'h0484: color = 2'b11;
      13'h0485: color = 2'b11;
      13'h0486: color = 2'b11;
      13'h0487: color = 2'b11;
      13'h0488: color = 2'b11;
      13'h0489: color = 2'b11;
      13'h048a: color = 2'b11;
      13'h048b: color = 2'b11;
      13'h048c: color = 2'b11;
      13'h048d: color = 2'b11;
      13'h048e: color = 2'b11;
      13'h048f: color = 2'b11;
      13'h0490: color = 2'b10;
      13'h0491: color = 2'b10;
      13'h0492: color = 2'b11;
      13'h0493: color = 2'b11;
      13'h0494: color = 2'b11;
      13'h0495: color = 2'b11;
      13'h0496: color = 2'b11;
      13'h0497: color = 2'b11;
      13'h0498: color = 2'b11;
      13'h0499: color = 2'b11;
      13'h049a: color = 2'b11;
      13'h049b: color = 2'b11;
      13'h049c: color = 2'b11;
      13'h049d: color = 2'b11;
      13'h049e: color = 2'b11;
      13'h049f: color = 2'b11;
      13'h04a0: color = 2'b00;
      13'h04a1: color = 2'b00;
      13'h04a2: color = 2'b11;
      13'h04a3: color = 2'b11;
      13'h04a4: color = 2'b10;
      13'h04a5: color = 2'b10;
      13'h04a6: color = 2'b10;
      13'h04a7: color = 2'b10;
      13'h04a8: color = 2'b10;
      13'h04a9: color = 2'b10;
      13'h04aa: color = 2'b10;
      13'h04ab: color = 2'b10;
      13'h04ac: color = 2'b10;
      13'h04ad: color = 2'b10;
      13'h04ae: color = 2'b10;
      13'h04af: color = 2'b10;
      13'h04b0: color = 2'b10;
      13'h04b1: color = 2'b10;
      13'h04b2: color = 2'b10;
      13'h04b3: color = 2'b10;
      13'h04b4: color = 2'b10;
      13'h04b5: color = 2'b10;
      13'h04b6: color = 2'b10;
      13'h04b7: color = 2'b10;
      13'h04b8: color = 2'b10;
      13'h04b9: color = 2'b10;
      13'h04ba: color = 2'b10;
      13'h04bb: color = 2'b10;
      13'h04bc: color = 2'b10;
      13'h04bd: color = 2'b10;
      13'h04be: color = 2'b10;
      13'h04bf: color = 2'b10;
      13'h04c0: color = 2'b10;
      13'h04c1: color = 2'b10;
      13'h04c2: color = 2'b10;
      13'h04c3: color = 2'b10;
      13'h04c4: color = 2'b10;
      13'h04c5: color = 2'b10;
      13'h04c6: color = 2'b10;
      13'h04c7: color = 2'b10;
      13'h04c8: color = 2'b10;
      13'h04c9: color = 2'b10;
      13'h04ca: color = 2'b10;
      13'h04cb: color = 2'b10;
      13'h04cc: color = 2'b10;
      13'h04cd: color = 2'b10;
      13'h04ce: color = 2'b10;
      13'h04cf: color = 2'b10;
      13'h04d0: color = 2'b10;
      13'h04d1: color = 2'b10;
      13'h04d2: color = 2'b10;
      13'h04d3: color = 2'b10;
      13'h04d4: color = 2'b10;
      13'h04d5: color = 2'b10;
      13'h04d6: color = 2'b10;
      13'h04d7: color = 2'b10;
      13'h04d8: color = 2'b10;
      13'h04d9: color = 2'b10;
      13'h04da: color = 2'b10;
      13'h04db: color = 2'b10;
      13'h04dc: color = 2'b01;
      13'h04dd: color = 2'b01;
      13'h04de: color = 2'b00;
      13'h04df: color = 2'b00;
      13'h04e0: color = 2'b10;
      13'h04e1: color = 2'b10;
      13'h04e2: color = 2'b11;
      13'h04e3: color = 2'b11;
      13'h04e4: color = 2'b11;
      13'h04e5: color = 2'b11;
      13'h04e6: color = 2'b11;
      13'h04e7: color = 2'b11;
      13'h04e8: color = 2'b11;
      13'h04e9: color = 2'b11;
      13'h04ea: color = 2'b11;
      13'h04eb: color = 2'b11;
      13'h04ec: color = 2'b11;
      13'h04ed: color = 2'b11;
      13'h04ee: color = 2'b11;
      13'h04ef: color = 2'b11;
      13'h04f0: color = 2'b10;
      13'h04f1: color = 2'b10;
      13'h04f2: color = 2'b11;
      13'h04f3: color = 2'b11;
      13'h04f4: color = 2'b11;
      13'h04f5: color = 2'b11;
      13'h04f6: color = 2'b11;
      13'h04f7: color = 2'b11;
      13'h04f8: color = 2'b11;
      13'h04f9: color = 2'b11;
      13'h04fa: color = 2'b11;
      13'h04fb: color = 2'b11;
      13'h04fc: color = 2'b11;
      13'h04fd: color = 2'b11;
      13'h04fe: color = 2'b11;
      13'h04ff: color = 2'b11;
      13'h0500: color = 2'b11;
      13'h0501: color = 2'b11;
      13'h0502: color = 2'b10;
      13'h0503: color = 2'b10;
      13'h0504: color = 2'b11;
      13'h0505: color = 2'b11;
      13'h0506: color = 2'b00;
      13'h0507: color = 2'b00;
      13'h0508: color = 2'b00;
      13'h0509: color = 2'b00;
      13'h050a: color = 2'b00;
      13'h050b: color = 2'b00;
      13'h050c: color = 2'b00;
      13'h050d: color = 2'b00;
      13'h050e: color = 2'b00;
      13'h050f: color = 2'b00;
      13'h0510: color = 2'b00;
      13'h0511: color = 2'b00;
      13'h0512: color = 2'b00;
      13'h0513: color = 2'b00;
      13'h0514: color = 2'b00;
      13'h0515: color = 2'b00;
      13'h0516: color = 2'b00;
      13'h0517: color = 2'b00;
      13'h0518: color = 2'b00;
      13'h0519: color = 2'b00;
      13'h051a: color = 2'b11;
      13'h051b: color = 2'b11;
      13'h051c: color = 2'b11;
      13'h051d: color = 2'b11;
      13'h051e: color = 2'b11;
      13'h051f: color = 2'b11;
      13'h0520: color = 2'b00;
      13'h0521: color = 2'b00;
      13'h0522: color = 2'b11;
      13'h0523: color = 2'b11;
      13'h0524: color = 2'b10;
      13'h0525: color = 2'b10;
      13'h0526: color = 2'b10;
      13'h0527: color = 2'b10;
      13'h0528: color = 2'b10;
      13'h0529: color = 2'b10;
      13'h052a: color = 2'b10;
      13'h052b: color = 2'b10;
      13'h052c: color = 2'b10;
      13'h052d: color = 2'b10;
      13'h052e: color = 2'b10;
      13'h052f: color = 2'b10;
      13'h0530: color = 2'b10;
      13'h0531: color = 2'b10;
      13'h0532: color = 2'b10;
      13'h0533: color = 2'b10;
      13'h0534: color = 2'b10;
      13'h0535: color = 2'b10;
      13'h0536: color = 2'b10;
      13'h0537: color = 2'b10;
      13'h0538: color = 2'b10;
      13'h0539: color = 2'b10;
      13'h053a: color = 2'b10;
      13'h053b: color = 2'b10;
      13'h053c: color = 2'b10;
      13'h053d: color = 2'b10;
      13'h053e: color = 2'b10;
      13'h053f: color = 2'b10;
      13'h0540: color = 2'b10;
      13'h0541: color = 2'b10;
      13'h0542: color = 2'b10;
      13'h0543: color = 2'b10;
      13'h0544: color = 2'b10;
      13'h0545: color = 2'b10;
      13'h0546: color = 2'b10;
      13'h0547: color = 2'b10;
      13'h0548: color = 2'b10;
      13'h0549: color = 2'b10;
      13'h054a: color = 2'b10;
      13'h054b: color = 2'b10;
      13'h054c: color = 2'b10;
      13'h054d: color = 2'b10;
      13'h054e: color = 2'b10;
      13'h054f: color = 2'b10;
      13'h0550: color = 2'b10;
      13'h0551: color = 2'b10;
      13'h0552: color = 2'b10;
      13'h0553: color = 2'b10;
      13'h0554: color = 2'b10;
      13'h0555: color = 2'b10;
      13'h0556: color = 2'b10;
      13'h0557: color = 2'b10;
      13'h0558: color = 2'b10;
      13'h0559: color = 2'b10;
      13'h055a: color = 2'b10;
      13'h055b: color = 2'b10;
      13'h055c: color = 2'b01;
      13'h055d: color = 2'b01;
      13'h055e: color = 2'b00;
      13'h055f: color = 2'b00;
      13'h0560: color = 2'b11;
      13'h0561: color = 2'b11;
      13'h0562: color = 2'b10;
      13'h0563: color = 2'b10;
      13'h0564: color = 2'b11;
      13'h0565: color = 2'b11;
      13'h0566: color = 2'b00;
      13'h0567: color = 2'b00;
      13'h0568: color = 2'b00;
      13'h0569: color = 2'b00;
      13'h056a: color = 2'b00;
      13'h056b: color = 2'b00;
      13'h056c: color = 2'b00;
      13'h056d: color = 2'b00;
      13'h056e: color = 2'b00;
      13'h056f: color = 2'b00;
      13'h0570: color = 2'b00;
      13'h0571: color = 2'b00;
      13'h0572: color = 2'b00;
      13'h0573: color = 2'b00;
      13'h0574: color = 2'b00;
      13'h0575: color = 2'b00;
      13'h0576: color = 2'b00;
      13'h0577: color = 2'b00;
      13'h0578: color = 2'b00;
      13'h0579: color = 2'b00;
      13'h057a: color = 2'b11;
      13'h057b: color = 2'b11;
      13'h057c: color = 2'b11;
      13'h057d: color = 2'b11;
      13'h057e: color = 2'b11;
      13'h057f: color = 2'b11;
      13'h0580: color = 2'b11;
      13'h0581: color = 2'b11;
      13'h0582: color = 2'b10;
      13'h0583: color = 2'b10;
      13'h0584: color = 2'b11;
      13'h0585: color = 2'b11;
      13'h0586: color = 2'b00;
      13'h0587: color = 2'b00;
      13'h0588: color = 2'b00;
      13'h0589: color = 2'b00;
      13'h058a: color = 2'b00;
      13'h058b: color = 2'b00;
      13'h058c: color = 2'b00;
      13'h058d: color = 2'b00;
      13'h058e: color = 2'b00;
      13'h058f: color = 2'b00;
      13'h0590: color = 2'b00;
      13'h0591: color = 2'b00;
      13'h0592: color = 2'b00;
      13'h0593: color = 2'b00;
      13'h0594: color = 2'b00;
      13'h0595: color = 2'b00;
      13'h0596: color = 2'b00;
      13'h0597: color = 2'b00;
      13'h0598: color = 2'b00;
      13'h0599: color = 2'b00;
      13'h059a: color = 2'b11;
      13'h059b: color = 2'b11;
      13'h059c: color = 2'b11;
      13'h059d: color = 2'b11;
      13'h059e: color = 2'b11;
      13'h059f: color = 2'b11;
      13'h05a0: color = 2'b00;
      13'h05a1: color = 2'b00;
      13'h05a2: color = 2'b11;
      13'h05a3: color = 2'b11;
      13'h05a4: color = 2'b10;
      13'h05a5: color = 2'b10;
      13'h05a6: color = 2'b10;
      13'h05a7: color = 2'b10;
      13'h05a8: color = 2'b10;
      13'h05a9: color = 2'b10;
      13'h05aa: color = 2'b10;
      13'h05ab: color = 2'b10;
      13'h05ac: color = 2'b10;
      13'h05ad: color = 2'b10;
      13'h05ae: color = 2'b10;
      13'h05af: color = 2'b10;
      13'h05b0: color = 2'b10;
      13'h05b1: color = 2'b10;
      13'h05b2: color = 2'b10;
      13'h05b3: color = 2'b10;
      13'h05b4: color = 2'b10;
      13'h05b5: color = 2'b10;
      13'h05b6: color = 2'b10;
      13'h05b7: color = 2'b10;
      13'h05b8: color = 2'b10;
      13'h05b9: color = 2'b10;
      13'h05ba: color = 2'b10;
      13'h05bb: color = 2'b10;
      13'h05bc: color = 2'b10;
      13'h05bd: color = 2'b10;
      13'h05be: color = 2'b10;
      13'h05bf: color = 2'b10;
      13'h05c0: color = 2'b10;
      13'h05c1: color = 2'b10;
      13'h05c2: color = 2'b10;
      13'h05c3: color = 2'b10;
      13'h05c4: color = 2'b10;
      13'h05c5: color = 2'b10;
      13'h05c6: color = 2'b10;
      13'h05c7: color = 2'b10;
      13'h05c8: color = 2'b10;
      13'h05c9: color = 2'b10;
      13'h05ca: color = 2'b10;
      13'h05cb: color = 2'b10;
      13'h05cc: color = 2'b10;
      13'h05cd: color = 2'b10;
      13'h05ce: color = 2'b10;
      13'h05cf: color = 2'b10;
      13'h05d0: color = 2'b10;
      13'h05d1: color = 2'b10;
      13'h05d2: color = 2'b10;
      13'h05d3: color = 2'b10;
      13'h05d4: color = 2'b10;
      13'h05d5: color = 2'b10;
      13'h05d6: color = 2'b10;
      13'h05d7: color = 2'b10;
      13'h05d8: color = 2'b10;
      13'h05d9: color = 2'b10;
      13'h05da: color = 2'b10;
      13'h05db: color = 2'b10;
      13'h05dc: color = 2'b01;
      13'h05dd: color = 2'b01;
      13'h05de: color = 2'b00;
      13'h05df: color = 2'b00;
      13'h05e0: color = 2'b11;
      13'h05e1: color = 2'b11;
      13'h05e2: color = 2'b10;
      13'h05e3: color = 2'b10;
      13'h05e4: color = 2'b11;
      13'h05e5: color = 2'b11;
      13'h05e6: color = 2'b00;
      13'h05e7: color = 2'b00;
      13'h05e8: color = 2'b00;
      13'h05e9: color = 2'b00;
      13'h05ea: color = 2'b00;
      13'h05eb: color = 2'b00;
      13'h05ec: color = 2'b00;
      13'h05ed: color = 2'b00;
      13'h05ee: color = 2'b00;
      13'h05ef: color = 2'b00;
      13'h05f0: color = 2'b00;
      13'h05f1: color = 2'b00;
      13'h05f2: color = 2'b00;
      13'h05f3: color = 2'b00;
      13'h05f4: color = 2'b00;
      13'h05f5: color = 2'b00;
      13'h05f6: color = 2'b00;
      13'h05f7: color = 2'b00;
      13'h05f8: color = 2'b00;
      13'h05f9: color = 2'b00;
      13'h05fa: color = 2'b11;
      13'h05fb: color = 2'b11;
      13'h05fc: color = 2'b11;
      13'h05fd: color = 2'b11;
      13'h05fe: color = 2'b11;
      13'h05ff: color = 2'b11;
      13'h0600: color = 2'b11;
      13'h0601: color = 2'b11;
      13'h0602: color = 2'b11;
      13'h0603: color = 2'b11;
      13'h0604: color = 2'b00;
      13'h0605: color = 2'b00;
      13'h0606: color = 2'b11;
      13'h0607: color = 2'b11;
      13'h0608: color = 2'b11;
      13'h0609: color = 2'b11;
      13'h060a: color = 2'b11;
      13'h060b: color = 2'b11;
      13'h060c: color = 2'b11;
      13'h060d: color = 2'b11;
      13'h060e: color = 2'b11;
      13'h060f: color = 2'b11;
      13'h0610: color = 2'b11;
      13'h0611: color = 2'b11;
      13'h0612: color = 2'b11;
      13'h0613: color = 2'b11;
      13'h0614: color = 2'b11;
      13'h0615: color = 2'b11;
      13'h0616: color = 2'b11;
      13'h0617: color = 2'b11;
      13'h0618: color = 2'b11;
      13'h0619: color = 2'b11;
      13'h061a: color = 2'b00;
      13'h061b: color = 2'b00;
      13'h061c: color = 2'b11;
      13'h061d: color = 2'b11;
      13'h061e: color = 2'b11;
      13'h061f: color = 2'b11;
      13'h0620: color = 2'b00;
      13'h0621: color = 2'b00;
      13'h0622: color = 2'b11;
      13'h0623: color = 2'b11;
      13'h0624: color = 2'b10;
      13'h0625: color = 2'b10;
      13'h0626: color = 2'b10;
      13'h0627: color = 2'b10;
      13'h0628: color = 2'b10;
      13'h0629: color = 2'b10;
      13'h062a: color = 2'b10;
      13'h062b: color = 2'b10;
      13'h062c: color = 2'b10;
      13'h062d: color = 2'b10;
      13'h062e: color = 2'b10;
      13'h062f: color = 2'b10;
      13'h0630: color = 2'b10;
      13'h0631: color = 2'b10;
      13'h0632: color = 2'b10;
      13'h0633: color = 2'b10;
      13'h0634: color = 2'b10;
      13'h0635: color = 2'b10;
      13'h0636: color = 2'b10;
      13'h0637: color = 2'b10;
      13'h0638: color = 2'b10;
      13'h0639: color = 2'b10;
      13'h063a: color = 2'b10;
      13'h063b: color = 2'b10;
      13'h063c: color = 2'b10;
      13'h063d: color = 2'b10;
      13'h063e: color = 2'b10;
      13'h063f: color = 2'b10;
      13'h0640: color = 2'b10;
      13'h0641: color = 2'b10;
      13'h0642: color = 2'b10;
      13'h0643: color = 2'b10;
      13'h0644: color = 2'b10;
      13'h0645: color = 2'b10;
      13'h0646: color = 2'b10;
      13'h0647: color = 2'b10;
      13'h0648: color = 2'b10;
      13'h0649: color = 2'b10;
      13'h064a: color = 2'b10;
      13'h064b: color = 2'b10;
      13'h064c: color = 2'b10;
      13'h064d: color = 2'b10;
      13'h064e: color = 2'b10;
      13'h064f: color = 2'b10;
      13'h0650: color = 2'b10;
      13'h0651: color = 2'b10;
      13'h0652: color = 2'b10;
      13'h0653: color = 2'b10;
      13'h0654: color = 2'b10;
      13'h0655: color = 2'b10;
      13'h0656: color = 2'b10;
      13'h0657: color = 2'b10;
      13'h0658: color = 2'b10;
      13'h0659: color = 2'b10;
      13'h065a: color = 2'b10;
      13'h065b: color = 2'b10;
      13'h065c: color = 2'b01;
      13'h065d: color = 2'b01;
      13'h065e: color = 2'b00;
      13'h065f: color = 2'b00;
      13'h0660: color = 2'b11;
      13'h0661: color = 2'b11;
      13'h0662: color = 2'b11;
      13'h0663: color = 2'b11;
      13'h0664: color = 2'b00;
      13'h0665: color = 2'b00;
      13'h0666: color = 2'b11;
      13'h0667: color = 2'b11;
      13'h0668: color = 2'b11;
      13'h0669: color = 2'b11;
      13'h066a: color = 2'b11;
      13'h066b: color = 2'b11;
      13'h066c: color = 2'b11;
      13'h066d: color = 2'b11;
      13'h066e: color = 2'b11;
      13'h066f: color = 2'b11;
      13'h0670: color = 2'b11;
      13'h0671: color = 2'b11;
      13'h0672: color = 2'b11;
      13'h0673: color = 2'b11;
      13'h0674: color = 2'b11;
      13'h0675: color = 2'b11;
      13'h0676: color = 2'b11;
      13'h0677: color = 2'b11;
      13'h0678: color = 2'b11;
      13'h0679: color = 2'b11;
      13'h067a: color = 2'b00;
      13'h067b: color = 2'b00;
      13'h067c: color = 2'b11;
      13'h067d: color = 2'b11;
      13'h067e: color = 2'b11;
      13'h067f: color = 2'b11;
      13'h0680: color = 2'b11;
      13'h0681: color = 2'b11;
      13'h0682: color = 2'b11;
      13'h0683: color = 2'b11;
      13'h0684: color = 2'b00;
      13'h0685: color = 2'b00;
      13'h0686: color = 2'b11;
      13'h0687: color = 2'b11;
      13'h0688: color = 2'b11;
      13'h0689: color = 2'b11;
      13'h068a: color = 2'b11;
      13'h068b: color = 2'b11;
      13'h068c: color = 2'b11;
      13'h068d: color = 2'b11;
      13'h068e: color = 2'b11;
      13'h068f: color = 2'b11;
      13'h0690: color = 2'b11;
      13'h0691: color = 2'b11;
      13'h0692: color = 2'b11;
      13'h0693: color = 2'b11;
      13'h0694: color = 2'b11;
      13'h0695: color = 2'b11;
      13'h0696: color = 2'b11;
      13'h0697: color = 2'b11;
      13'h0698: color = 2'b11;
      13'h0699: color = 2'b11;
      13'h069a: color = 2'b00;
      13'h069b: color = 2'b00;
      13'h069c: color = 2'b11;
      13'h069d: color = 2'b11;
      13'h069e: color = 2'b11;
      13'h069f: color = 2'b11;
      13'h06a0: color = 2'b00;
      13'h06a1: color = 2'b00;
      13'h06a2: color = 2'b11;
      13'h06a3: color = 2'b11;
      13'h06a4: color = 2'b10;
      13'h06a5: color = 2'b10;
      13'h06a6: color = 2'b10;
      13'h06a7: color = 2'b10;
      13'h06a8: color = 2'b10;
      13'h06a9: color = 2'b10;
      13'h06aa: color = 2'b10;
      13'h06ab: color = 2'b10;
      13'h06ac: color = 2'b10;
      13'h06ad: color = 2'b10;
      13'h06ae: color = 2'b10;
      13'h06af: color = 2'b10;
      13'h06b0: color = 2'b10;
      13'h06b1: color = 2'b10;
      13'h06b2: color = 2'b10;
      13'h06b3: color = 2'b10;
      13'h06b4: color = 2'b10;
      13'h06b5: color = 2'b10;
      13'h06b6: color = 2'b10;
      13'h06b7: color = 2'b10;
      13'h06b8: color = 2'b10;
      13'h06b9: color = 2'b10;
      13'h06ba: color = 2'b10;
      13'h06bb: color = 2'b10;
      13'h06bc: color = 2'b10;
      13'h06bd: color = 2'b10;
      13'h06be: color = 2'b10;
      13'h06bf: color = 2'b10;
      13'h06c0: color = 2'b10;
      13'h06c1: color = 2'b10;
      13'h06c2: color = 2'b10;
      13'h06c3: color = 2'b10;
      13'h06c4: color = 2'b10;
      13'h06c5: color = 2'b10;
      13'h06c6: color = 2'b10;
      13'h06c7: color = 2'b10;
      13'h06c8: color = 2'b10;
      13'h06c9: color = 2'b10;
      13'h06ca: color = 2'b10;
      13'h06cb: color = 2'b10;
      13'h06cc: color = 2'b10;
      13'h06cd: color = 2'b10;
      13'h06ce: color = 2'b10;
      13'h06cf: color = 2'b10;
      13'h06d0: color = 2'b10;
      13'h06d1: color = 2'b10;
      13'h06d2: color = 2'b10;
      13'h06d3: color = 2'b10;
      13'h06d4: color = 2'b10;
      13'h06d5: color = 2'b10;
      13'h06d6: color = 2'b10;
      13'h06d7: color = 2'b10;
      13'h06d8: color = 2'b10;
      13'h06d9: color = 2'b10;
      13'h06da: color = 2'b10;
      13'h06db: color = 2'b10;
      13'h06dc: color = 2'b01;
      13'h06dd: color = 2'b01;
      13'h06de: color = 2'b00;
      13'h06df: color = 2'b00;
      13'h06e0: color = 2'b11;
      13'h06e1: color = 2'b11;
      13'h06e2: color = 2'b11;
      13'h06e3: color = 2'b11;
      13'h06e4: color = 2'b00;
      13'h06e5: color = 2'b00;
      13'h06e6: color = 2'b11;
      13'h06e7: color = 2'b11;
      13'h06e8: color = 2'b11;
      13'h06e9: color = 2'b11;
      13'h06ea: color = 2'b11;
      13'h06eb: color = 2'b11;
      13'h06ec: color = 2'b11;
      13'h06ed: color = 2'b11;
      13'h06ee: color = 2'b11;
      13'h06ef: color = 2'b11;
      13'h06f0: color = 2'b11;
      13'h06f1: color = 2'b11;
      13'h06f2: color = 2'b11;
      13'h06f3: color = 2'b11;
      13'h06f4: color = 2'b11;
      13'h06f5: color = 2'b11;
      13'h06f6: color = 2'b11;
      13'h06f7: color = 2'b11;
      13'h06f8: color = 2'b11;
      13'h06f9: color = 2'b11;
      13'h06fa: color = 2'b00;
      13'h06fb: color = 2'b00;
      13'h06fc: color = 2'b11;
      13'h06fd: color = 2'b11;
      13'h06fe: color = 2'b11;
      13'h06ff: color = 2'b11;
      13'h0700: color = 2'b11;
      13'h0701: color = 2'b11;
      13'h0702: color = 2'b11;
      13'h0703: color = 2'b11;
      13'h0704: color = 2'b00;
      13'h0705: color = 2'b00;
      13'h0706: color = 2'b11;
      13'h0707: color = 2'b11;
      13'h0708: color = 2'b11;
      13'h0709: color = 2'b11;
      13'h070a: color = 2'b10;
      13'h070b: color = 2'b10;
      13'h070c: color = 2'b10;
      13'h070d: color = 2'b10;
      13'h070e: color = 2'b10;
      13'h070f: color = 2'b10;
      13'h0710: color = 2'b10;
      13'h0711: color = 2'b10;
      13'h0712: color = 2'b10;
      13'h0713: color = 2'b10;
      13'h0714: color = 2'b10;
      13'h0715: color = 2'b10;
      13'h0716: color = 2'b11;
      13'h0717: color = 2'b11;
      13'h0718: color = 2'b11;
      13'h0719: color = 2'b11;
      13'h071a: color = 2'b00;
      13'h071b: color = 2'b00;
      13'h071c: color = 2'b11;
      13'h071d: color = 2'b11;
      13'h071e: color = 2'b11;
      13'h071f: color = 2'b11;
      13'h0720: color = 2'b00;
      13'h0721: color = 2'b00;
      13'h0722: color = 2'b11;
      13'h0723: color = 2'b11;
      13'h0724: color = 2'b10;
      13'h0725: color = 2'b10;
      13'h0726: color = 2'b10;
      13'h0727: color = 2'b10;
      13'h0728: color = 2'b10;
      13'h0729: color = 2'b10;
      13'h072a: color = 2'b10;
      13'h072b: color = 2'b10;
      13'h072c: color = 2'b10;
      13'h072d: color = 2'b10;
      13'h072e: color = 2'b10;
      13'h072f: color = 2'b10;
      13'h0730: color = 2'b10;
      13'h0731: color = 2'b10;
      13'h0732: color = 2'b10;
      13'h0733: color = 2'b10;
      13'h0734: color = 2'b10;
      13'h0735: color = 2'b10;
      13'h0736: color = 2'b10;
      13'h0737: color = 2'b10;
      13'h0738: color = 2'b10;
      13'h0739: color = 2'b10;
      13'h073a: color = 2'b10;
      13'h073b: color = 2'b10;
      13'h073c: color = 2'b10;
      13'h073d: color = 2'b10;
      13'h073e: color = 2'b10;
      13'h073f: color = 2'b10;
      13'h0740: color = 2'b10;
      13'h0741: color = 2'b10;
      13'h0742: color = 2'b10;
      13'h0743: color = 2'b10;
      13'h0744: color = 2'b10;
      13'h0745: color = 2'b10;
      13'h0746: color = 2'b10;
      13'h0747: color = 2'b10;
      13'h0748: color = 2'b10;
      13'h0749: color = 2'b10;
      13'h074a: color = 2'b10;
      13'h074b: color = 2'b10;
      13'h074c: color = 2'b10;
      13'h074d: color = 2'b10;
      13'h074e: color = 2'b10;
      13'h074f: color = 2'b10;
      13'h0750: color = 2'b10;
      13'h0751: color = 2'b10;
      13'h0752: color = 2'b10;
      13'h0753: color = 2'b10;
      13'h0754: color = 2'b10;
      13'h0755: color = 2'b10;
      13'h0756: color = 2'b10;
      13'h0757: color = 2'b10;
      13'h0758: color = 2'b10;
      13'h0759: color = 2'b10;
      13'h075a: color = 2'b10;
      13'h075b: color = 2'b10;
      13'h075c: color = 2'b01;
      13'h075d: color = 2'b01;
      13'h075e: color = 2'b00;
      13'h075f: color = 2'b00;
      13'h0760: color = 2'b11;
      13'h0761: color = 2'b11;
      13'h0762: color = 2'b11;
      13'h0763: color = 2'b11;
      13'h0764: color = 2'b00;
      13'h0765: color = 2'b00;
      13'h0766: color = 2'b11;
      13'h0767: color = 2'b11;
      13'h0768: color = 2'b11;
      13'h0769: color = 2'b11;
      13'h076a: color = 2'b10;
      13'h076b: color = 2'b10;
      13'h076c: color = 2'b10;
      13'h076d: color = 2'b10;
      13'h076e: color = 2'b10;
      13'h076f: color = 2'b10;
      13'h0770: color = 2'b10;
      13'h0771: color = 2'b10;
      13'h0772: color = 2'b10;
      13'h0773: color = 2'b10;
      13'h0774: color = 2'b10;
      13'h0775: color = 2'b10;
      13'h0776: color = 2'b11;
      13'h0777: color = 2'b11;
      13'h0778: color = 2'b11;
      13'h0779: color = 2'b11;
      13'h077a: color = 2'b00;
      13'h077b: color = 2'b00;
      13'h077c: color = 2'b11;
      13'h077d: color = 2'b11;
      13'h077e: color = 2'b11;
      13'h077f: color = 2'b11;
      13'h0780: color = 2'b11;
      13'h0781: color = 2'b11;
      13'h0782: color = 2'b11;
      13'h0783: color = 2'b11;
      13'h0784: color = 2'b00;
      13'h0785: color = 2'b00;
      13'h0786: color = 2'b11;
      13'h0787: color = 2'b11;
      13'h0788: color = 2'b11;
      13'h0789: color = 2'b11;
      13'h078a: color = 2'b10;
      13'h078b: color = 2'b10;
      13'h078c: color = 2'b10;
      13'h078d: color = 2'b10;
      13'h078e: color = 2'b10;
      13'h078f: color = 2'b10;
      13'h0790: color = 2'b10;
      13'h0791: color = 2'b10;
      13'h0792: color = 2'b10;
      13'h0793: color = 2'b10;
      13'h0794: color = 2'b10;
      13'h0795: color = 2'b10;
      13'h0796: color = 2'b11;
      13'h0797: color = 2'b11;
      13'h0798: color = 2'b11;
      13'h0799: color = 2'b11;
      13'h079a: color = 2'b00;
      13'h079b: color = 2'b00;
      13'h079c: color = 2'b11;
      13'h079d: color = 2'b11;
      13'h079e: color = 2'b11;
      13'h079f: color = 2'b11;
      13'h07a0: color = 2'b00;
      13'h07a1: color = 2'b00;
      13'h07a2: color = 2'b11;
      13'h07a3: color = 2'b11;
      13'h07a4: color = 2'b10;
      13'h07a5: color = 2'b10;
      13'h07a6: color = 2'b10;
      13'h07a7: color = 2'b10;
      13'h07a8: color = 2'b10;
      13'h07a9: color = 2'b10;
      13'h07aa: color = 2'b10;
      13'h07ab: color = 2'b10;
      13'h07ac: color = 2'b10;
      13'h07ad: color = 2'b10;
      13'h07ae: color = 2'b10;
      13'h07af: color = 2'b10;
      13'h07b0: color = 2'b10;
      13'h07b1: color = 2'b10;
      13'h07b2: color = 2'b10;
      13'h07b3: color = 2'b10;
      13'h07b4: color = 2'b10;
      13'h07b5: color = 2'b10;
      13'h07b6: color = 2'b10;
      13'h07b7: color = 2'b10;
      13'h07b8: color = 2'b10;
      13'h07b9: color = 2'b10;
      13'h07ba: color = 2'b10;
      13'h07bb: color = 2'b10;
      13'h07bc: color = 2'b10;
      13'h07bd: color = 2'b10;
      13'h07be: color = 2'b10;
      13'h07bf: color = 2'b10;
      13'h07c0: color = 2'b10;
      13'h07c1: color = 2'b10;
      13'h07c2: color = 2'b10;
      13'h07c3: color = 2'b10;
      13'h07c4: color = 2'b10;
      13'h07c5: color = 2'b10;
      13'h07c6: color = 2'b10;
      13'h07c7: color = 2'b10;
      13'h07c8: color = 2'b10;
      13'h07c9: color = 2'b10;
      13'h07ca: color = 2'b10;
      13'h07cb: color = 2'b10;
      13'h07cc: color = 2'b10;
      13'h07cd: color = 2'b10;
      13'h07ce: color = 2'b10;
      13'h07cf: color = 2'b10;
      13'h07d0: color = 2'b10;
      13'h07d1: color = 2'b10;
      13'h07d2: color = 2'b10;
      13'h07d3: color = 2'b10;
      13'h07d4: color = 2'b10;
      13'h07d5: color = 2'b10;
      13'h07d6: color = 2'b10;
      13'h07d7: color = 2'b10;
      13'h07d8: color = 2'b10;
      13'h07d9: color = 2'b10;
      13'h07da: color = 2'b10;
      13'h07db: color = 2'b10;
      13'h07dc: color = 2'b01;
      13'h07dd: color = 2'b01;
      13'h07de: color = 2'b00;
      13'h07df: color = 2'b00;
      13'h07e0: color = 2'b11;
      13'h07e1: color = 2'b11;
      13'h07e2: color = 2'b11;
      13'h07e3: color = 2'b11;
      13'h07e4: color = 2'b00;
      13'h07e5: color = 2'b00;
      13'h07e6: color = 2'b11;
      13'h07e7: color = 2'b11;
      13'h07e8: color = 2'b11;
      13'h07e9: color = 2'b11;
      13'h07ea: color = 2'b10;
      13'h07eb: color = 2'b10;
      13'h07ec: color = 2'b10;
      13'h07ed: color = 2'b10;
      13'h07ee: color = 2'b10;
      13'h07ef: color = 2'b10;
      13'h07f0: color = 2'b10;
      13'h07f1: color = 2'b10;
      13'h07f2: color = 2'b10;
      13'h07f3: color = 2'b10;
      13'h07f4: color = 2'b10;
      13'h07f5: color = 2'b10;
      13'h07f6: color = 2'b11;
      13'h07f7: color = 2'b11;
      13'h07f8: color = 2'b11;
      13'h07f9: color = 2'b11;
      13'h07fa: color = 2'b00;
      13'h07fb: color = 2'b00;
      13'h07fc: color = 2'b11;
      13'h07fd: color = 2'b11;
      13'h07fe: color = 2'b11;
      13'h07ff: color = 2'b11;
      13'h0800: color = 2'b11;
      13'h0801: color = 2'b11;
      13'h0802: color = 2'b11;
      13'h0803: color = 2'b11;
      13'h0804: color = 2'b00;
      13'h0805: color = 2'b00;
      13'h0806: color = 2'b11;
      13'h0807: color = 2'b11;
      13'h0808: color = 2'b11;
      13'h0809: color = 2'b11;
      13'h080a: color = 2'b10;
      13'h080b: color = 2'b10;
      13'h080c: color = 2'b10;
      13'h080d: color = 2'b10;
      13'h080e: color = 2'b10;
      13'h080f: color = 2'b10;
      13'h0810: color = 2'b10;
      13'h0811: color = 2'b10;
      13'h0812: color = 2'b10;
      13'h0813: color = 2'b10;
      13'h0814: color = 2'b10;
      13'h0815: color = 2'b10;
      13'h0816: color = 2'b11;
      13'h0817: color = 2'b11;
      13'h0818: color = 2'b11;
      13'h0819: color = 2'b11;
      13'h081a: color = 2'b00;
      13'h081b: color = 2'b00;
      13'h081c: color = 2'b11;
      13'h081d: color = 2'b11;
      13'h081e: color = 2'b11;
      13'h081f: color = 2'b11;
      13'h0820: color = 2'b00;
      13'h0821: color = 2'b00;
      13'h0822: color = 2'b11;
      13'h0823: color = 2'b11;
      13'h0824: color = 2'b10;
      13'h0825: color = 2'b10;
      13'h0826: color = 2'b10;
      13'h0827: color = 2'b10;
      13'h0828: color = 2'b10;
      13'h0829: color = 2'b10;
      13'h082a: color = 2'b10;
      13'h082b: color = 2'b10;
      13'h082c: color = 2'b10;
      13'h082d: color = 2'b10;
      13'h082e: color = 2'b10;
      13'h082f: color = 2'b10;
      13'h0830: color = 2'b10;
      13'h0831: color = 2'b10;
      13'h0832: color = 2'b10;
      13'h0833: color = 2'b10;
      13'h0834: color = 2'b10;
      13'h0835: color = 2'b10;
      13'h0836: color = 2'b10;
      13'h0837: color = 2'b10;
      13'h0838: color = 2'b10;
      13'h0839: color = 2'b10;
      13'h083a: color = 2'b10;
      13'h083b: color = 2'b10;
      13'h083c: color = 2'b10;
      13'h083d: color = 2'b10;
      13'h083e: color = 2'b10;
      13'h083f: color = 2'b10;
      13'h0840: color = 2'b10;
      13'h0841: color = 2'b10;
      13'h0842: color = 2'b10;
      13'h0843: color = 2'b10;
      13'h0844: color = 2'b10;
      13'h0845: color = 2'b10;
      13'h0846: color = 2'b10;
      13'h0847: color = 2'b10;
      13'h0848: color = 2'b10;
      13'h0849: color = 2'b10;
      13'h084a: color = 2'b10;
      13'h084b: color = 2'b10;
      13'h084c: color = 2'b10;
      13'h084d: color = 2'b10;
      13'h084e: color = 2'b10;
      13'h084f: color = 2'b10;
      13'h0850: color = 2'b10;
      13'h0851: color = 2'b10;
      13'h0852: color = 2'b10;
      13'h0853: color = 2'b10;
      13'h0854: color = 2'b10;
      13'h0855: color = 2'b10;
      13'h0856: color = 2'b10;
      13'h0857: color = 2'b10;
      13'h0858: color = 2'b10;
      13'h0859: color = 2'b10;
      13'h085a: color = 2'b10;
      13'h085b: color = 2'b10;
      13'h085c: color = 2'b01;
      13'h085d: color = 2'b01;
      13'h085e: color = 2'b00;
      13'h085f: color = 2'b00;
      13'h0860: color = 2'b11;
      13'h0861: color = 2'b11;
      13'h0862: color = 2'b11;
      13'h0863: color = 2'b11;
      13'h0864: color = 2'b00;
      13'h0865: color = 2'b00;
      13'h0866: color = 2'b11;
      13'h0867: color = 2'b11;
      13'h0868: color = 2'b11;
      13'h0869: color = 2'b11;
      13'h086a: color = 2'b10;
      13'h086b: color = 2'b10;
      13'h086c: color = 2'b10;
      13'h086d: color = 2'b10;
      13'h086e: color = 2'b10;
      13'h086f: color = 2'b10;
      13'h0870: color = 2'b10;
      13'h0871: color = 2'b10;
      13'h0872: color = 2'b10;
      13'h0873: color = 2'b10;
      13'h0874: color = 2'b10;
      13'h0875: color = 2'b10;
      13'h0876: color = 2'b11;
      13'h0877: color = 2'b11;
      13'h0878: color = 2'b11;
      13'h0879: color = 2'b11;
      13'h087a: color = 2'b00;
      13'h087b: color = 2'b00;
      13'h087c: color = 2'b11;
      13'h087d: color = 2'b11;
      13'h087e: color = 2'b11;
      13'h087f: color = 2'b11;
      13'h0880: color = 2'b11;
      13'h0881: color = 2'b11;
      13'h0882: color = 2'b11;
      13'h0883: color = 2'b11;
      13'h0884: color = 2'b00;
      13'h0885: color = 2'b00;
      13'h0886: color = 2'b11;
      13'h0887: color = 2'b11;
      13'h0888: color = 2'b11;
      13'h0889: color = 2'b11;
      13'h088a: color = 2'b10;
      13'h088b: color = 2'b10;
      13'h088c: color = 2'b10;
      13'h088d: color = 2'b10;
      13'h088e: color = 2'b10;
      13'h088f: color = 2'b10;
      13'h0890: color = 2'b10;
      13'h0891: color = 2'b10;
      13'h0892: color = 2'b10;
      13'h0893: color = 2'b10;
      13'h0894: color = 2'b10;
      13'h0895: color = 2'b10;
      13'h0896: color = 2'b11;
      13'h0897: color = 2'b11;
      13'h0898: color = 2'b11;
      13'h0899: color = 2'b11;
      13'h089a: color = 2'b00;
      13'h089b: color = 2'b00;
      13'h089c: color = 2'b11;
      13'h089d: color = 2'b11;
      13'h089e: color = 2'b11;
      13'h089f: color = 2'b11;
      13'h08a0: color = 2'b00;
      13'h08a1: color = 2'b00;
      13'h08a2: color = 2'b11;
      13'h08a3: color = 2'b11;
      13'h08a4: color = 2'b10;
      13'h08a5: color = 2'b10;
      13'h08a6: color = 2'b10;
      13'h08a7: color = 2'b10;
      13'h08a8: color = 2'b10;
      13'h08a9: color = 2'b10;
      13'h08aa: color = 2'b10;
      13'h08ab: color = 2'b10;
      13'h08ac: color = 2'b10;
      13'h08ad: color = 2'b10;
      13'h08ae: color = 2'b10;
      13'h08af: color = 2'b10;
      13'h08b0: color = 2'b10;
      13'h08b1: color = 2'b10;
      13'h08b2: color = 2'b10;
      13'h08b3: color = 2'b10;
      13'h08b4: color = 2'b10;
      13'h08b5: color = 2'b10;
      13'h08b6: color = 2'b10;
      13'h08b7: color = 2'b10;
      13'h08b8: color = 2'b10;
      13'h08b9: color = 2'b10;
      13'h08ba: color = 2'b10;
      13'h08bb: color = 2'b10;
      13'h08bc: color = 2'b10;
      13'h08bd: color = 2'b10;
      13'h08be: color = 2'b10;
      13'h08bf: color = 2'b10;
      13'h08c0: color = 2'b10;
      13'h08c1: color = 2'b10;
      13'h08c2: color = 2'b10;
      13'h08c3: color = 2'b10;
      13'h08c4: color = 2'b10;
      13'h08c5: color = 2'b10;
      13'h08c6: color = 2'b10;
      13'h08c7: color = 2'b10;
      13'h08c8: color = 2'b10;
      13'h08c9: color = 2'b10;
      13'h08ca: color = 2'b10;
      13'h08cb: color = 2'b10;
      13'h08cc: color = 2'b10;
      13'h08cd: color = 2'b10;
      13'h08ce: color = 2'b10;
      13'h08cf: color = 2'b10;
      13'h08d0: color = 2'b10;
      13'h08d1: color = 2'b10;
      13'h08d2: color = 2'b10;
      13'h08d3: color = 2'b10;
      13'h08d4: color = 2'b10;
      13'h08d5: color = 2'b10;
      13'h08d6: color = 2'b10;
      13'h08d7: color = 2'b10;
      13'h08d8: color = 2'b10;
      13'h08d9: color = 2'b10;
      13'h08da: color = 2'b10;
      13'h08db: color = 2'b10;
      13'h08dc: color = 2'b01;
      13'h08dd: color = 2'b01;
      13'h08de: color = 2'b00;
      13'h08df: color = 2'b00;
      13'h08e0: color = 2'b11;
      13'h08e1: color = 2'b11;
      13'h08e2: color = 2'b11;
      13'h08e3: color = 2'b11;
      13'h08e4: color = 2'b00;
      13'h08e5: color = 2'b00;
      13'h08e6: color = 2'b11;
      13'h08e7: color = 2'b11;
      13'h08e8: color = 2'b11;
      13'h08e9: color = 2'b11;
      13'h08ea: color = 2'b10;
      13'h08eb: color = 2'b10;
      13'h08ec: color = 2'b10;
      13'h08ed: color = 2'b10;
      13'h08ee: color = 2'b10;
      13'h08ef: color = 2'b10;
      13'h08f0: color = 2'b10;
      13'h08f1: color = 2'b10;
      13'h08f2: color = 2'b10;
      13'h08f3: color = 2'b10;
      13'h08f4: color = 2'b10;
      13'h08f5: color = 2'b10;
      13'h08f6: color = 2'b11;
      13'h08f7: color = 2'b11;
      13'h08f8: color = 2'b11;
      13'h08f9: color = 2'b11;
      13'h08fa: color = 2'b00;
      13'h08fb: color = 2'b00;
      13'h08fc: color = 2'b11;
      13'h08fd: color = 2'b11;
      13'h08fe: color = 2'b11;
      13'h08ff: color = 2'b11;
      13'h0900: color = 2'b11;
      13'h0901: color = 2'b11;
      13'h0902: color = 2'b10;
      13'h0903: color = 2'b10;
      13'h0904: color = 2'b00;
      13'h0905: color = 2'b00;
      13'h0906: color = 2'b11;
      13'h0907: color = 2'b11;
      13'h0908: color = 2'b11;
      13'h0909: color = 2'b11;
      13'h090a: color = 2'b10;
      13'h090b: color = 2'b10;
      13'h090c: color = 2'b10;
      13'h090d: color = 2'b10;
      13'h090e: color = 2'b10;
      13'h090f: color = 2'b10;
      13'h0910: color = 2'b10;
      13'h0911: color = 2'b10;
      13'h0912: color = 2'b10;
      13'h0913: color = 2'b10;
      13'h0914: color = 2'b10;
      13'h0915: color = 2'b10;
      13'h0916: color = 2'b11;
      13'h0917: color = 2'b11;
      13'h0918: color = 2'b11;
      13'h0919: color = 2'b11;
      13'h091a: color = 2'b00;
      13'h091b: color = 2'b00;
      13'h091c: color = 2'b11;
      13'h091d: color = 2'b11;
      13'h091e: color = 2'b11;
      13'h091f: color = 2'b11;
      13'h0920: color = 2'b00;
      13'h0921: color = 2'b00;
      13'h0922: color = 2'b11;
      13'h0923: color = 2'b11;
      13'h0924: color = 2'b10;
      13'h0925: color = 2'b10;
      13'h0926: color = 2'b10;
      13'h0927: color = 2'b10;
      13'h0928: color = 2'b10;
      13'h0929: color = 2'b10;
      13'h092a: color = 2'b10;
      13'h092b: color = 2'b10;
      13'h092c: color = 2'b10;
      13'h092d: color = 2'b10;
      13'h092e: color = 2'b10;
      13'h092f: color = 2'b10;
      13'h0930: color = 2'b10;
      13'h0931: color = 2'b10;
      13'h0932: color = 2'b10;
      13'h0933: color = 2'b10;
      13'h0934: color = 2'b10;
      13'h0935: color = 2'b10;
      13'h0936: color = 2'b10;
      13'h0937: color = 2'b10;
      13'h0938: color = 2'b10;
      13'h0939: color = 2'b10;
      13'h093a: color = 2'b10;
      13'h093b: color = 2'b10;
      13'h093c: color = 2'b10;
      13'h093d: color = 2'b10;
      13'h093e: color = 2'b10;
      13'h093f: color = 2'b10;
      13'h0940: color = 2'b10;
      13'h0941: color = 2'b10;
      13'h0942: color = 2'b10;
      13'h0943: color = 2'b10;
      13'h0944: color = 2'b10;
      13'h0945: color = 2'b10;
      13'h0946: color = 2'b10;
      13'h0947: color = 2'b10;
      13'h0948: color = 2'b10;
      13'h0949: color = 2'b10;
      13'h094a: color = 2'b10;
      13'h094b: color = 2'b10;
      13'h094c: color = 2'b10;
      13'h094d: color = 2'b10;
      13'h094e: color = 2'b10;
      13'h094f: color = 2'b10;
      13'h0950: color = 2'b10;
      13'h0951: color = 2'b10;
      13'h0952: color = 2'b10;
      13'h0953: color = 2'b10;
      13'h0954: color = 2'b10;
      13'h0955: color = 2'b10;
      13'h0956: color = 2'b10;
      13'h0957: color = 2'b10;
      13'h0958: color = 2'b10;
      13'h0959: color = 2'b10;
      13'h095a: color = 2'b10;
      13'h095b: color = 2'b10;
      13'h095c: color = 2'b01;
      13'h095d: color = 2'b01;
      13'h095e: color = 2'b00;
      13'h095f: color = 2'b00;
      13'h0960: color = 2'b11;
      13'h0961: color = 2'b11;
      13'h0962: color = 2'b10;
      13'h0963: color = 2'b10;
      13'h0964: color = 2'b00;
      13'h0965: color = 2'b00;
      13'h0966: color = 2'b11;
      13'h0967: color = 2'b11;
      13'h0968: color = 2'b11;
      13'h0969: color = 2'b11;
      13'h096a: color = 2'b10;
      13'h096b: color = 2'b10;
      13'h096c: color = 2'b10;
      13'h096d: color = 2'b10;
      13'h096e: color = 2'b10;
      13'h096f: color = 2'b10;
      13'h0970: color = 2'b10;
      13'h0971: color = 2'b10;
      13'h0972: color = 2'b10;
      13'h0973: color = 2'b10;
      13'h0974: color = 2'b10;
      13'h0975: color = 2'b10;
      13'h0976: color = 2'b11;
      13'h0977: color = 2'b11;
      13'h0978: color = 2'b11;
      13'h0979: color = 2'b11;
      13'h097a: color = 2'b00;
      13'h097b: color = 2'b00;
      13'h097c: color = 2'b11;
      13'h097d: color = 2'b11;
      13'h097e: color = 2'b11;
      13'h097f: color = 2'b11;
      13'h0980: color = 2'b11;
      13'h0981: color = 2'b11;
      13'h0982: color = 2'b10;
      13'h0983: color = 2'b10;
      13'h0984: color = 2'b00;
      13'h0985: color = 2'b00;
      13'h0986: color = 2'b11;
      13'h0987: color = 2'b11;
      13'h0988: color = 2'b11;
      13'h0989: color = 2'b11;
      13'h098a: color = 2'b10;
      13'h098b: color = 2'b10;
      13'h098c: color = 2'b10;
      13'h098d: color = 2'b10;
      13'h098e: color = 2'b10;
      13'h098f: color = 2'b10;
      13'h0990: color = 2'b10;
      13'h0991: color = 2'b10;
      13'h0992: color = 2'b10;
      13'h0993: color = 2'b10;
      13'h0994: color = 2'b10;
      13'h0995: color = 2'b10;
      13'h0996: color = 2'b11;
      13'h0997: color = 2'b11;
      13'h0998: color = 2'b11;
      13'h0999: color = 2'b11;
      13'h099a: color = 2'b00;
      13'h099b: color = 2'b00;
      13'h099c: color = 2'b11;
      13'h099d: color = 2'b11;
      13'h099e: color = 2'b11;
      13'h099f: color = 2'b11;
      13'h09a0: color = 2'b00;
      13'h09a1: color = 2'b00;
      13'h09a2: color = 2'b11;
      13'h09a3: color = 2'b11;
      13'h09a4: color = 2'b10;
      13'h09a5: color = 2'b10;
      13'h09a6: color = 2'b10;
      13'h09a7: color = 2'b10;
      13'h09a8: color = 2'b10;
      13'h09a9: color = 2'b10;
      13'h09aa: color = 2'b10;
      13'h09ab: color = 2'b10;
      13'h09ac: color = 2'b10;
      13'h09ad: color = 2'b10;
      13'h09ae: color = 2'b10;
      13'h09af: color = 2'b10;
      13'h09b0: color = 2'b10;
      13'h09b1: color = 2'b10;
      13'h09b2: color = 2'b10;
      13'h09b3: color = 2'b10;
      13'h09b4: color = 2'b10;
      13'h09b5: color = 2'b10;
      13'h09b6: color = 2'b10;
      13'h09b7: color = 2'b10;
      13'h09b8: color = 2'b10;
      13'h09b9: color = 2'b10;
      13'h09ba: color = 2'b10;
      13'h09bb: color = 2'b10;
      13'h09bc: color = 2'b10;
      13'h09bd: color = 2'b10;
      13'h09be: color = 2'b10;
      13'h09bf: color = 2'b10;
      13'h09c0: color = 2'b10;
      13'h09c1: color = 2'b10;
      13'h09c2: color = 2'b10;
      13'h09c3: color = 2'b10;
      13'h09c4: color = 2'b10;
      13'h09c5: color = 2'b10;
      13'h09c6: color = 2'b10;
      13'h09c7: color = 2'b10;
      13'h09c8: color = 2'b10;
      13'h09c9: color = 2'b10;
      13'h09ca: color = 2'b10;
      13'h09cb: color = 2'b10;
      13'h09cc: color = 2'b10;
      13'h09cd: color = 2'b10;
      13'h09ce: color = 2'b10;
      13'h09cf: color = 2'b10;
      13'h09d0: color = 2'b10;
      13'h09d1: color = 2'b10;
      13'h09d2: color = 2'b10;
      13'h09d3: color = 2'b10;
      13'h09d4: color = 2'b10;
      13'h09d5: color = 2'b10;
      13'h09d6: color = 2'b10;
      13'h09d7: color = 2'b10;
      13'h09d8: color = 2'b10;
      13'h09d9: color = 2'b10;
      13'h09da: color = 2'b10;
      13'h09db: color = 2'b10;
      13'h09dc: color = 2'b01;
      13'h09dd: color = 2'b01;
      13'h09de: color = 2'b00;
      13'h09df: color = 2'b00;
      13'h09e0: color = 2'b11;
      13'h09e1: color = 2'b11;
      13'h09e2: color = 2'b10;
      13'h09e3: color = 2'b10;
      13'h09e4: color = 2'b00;
      13'h09e5: color = 2'b00;
      13'h09e6: color = 2'b11;
      13'h09e7: color = 2'b11;
      13'h09e8: color = 2'b11;
      13'h09e9: color = 2'b11;
      13'h09ea: color = 2'b10;
      13'h09eb: color = 2'b10;
      13'h09ec: color = 2'b10;
      13'h09ed: color = 2'b10;
      13'h09ee: color = 2'b10;
      13'h09ef: color = 2'b10;
      13'h09f0: color = 2'b10;
      13'h09f1: color = 2'b10;
      13'h09f2: color = 2'b10;
      13'h09f3: color = 2'b10;
      13'h09f4: color = 2'b10;
      13'h09f5: color = 2'b10;
      13'h09f6: color = 2'b11;
      13'h09f7: color = 2'b11;
      13'h09f8: color = 2'b11;
      13'h09f9: color = 2'b11;
      13'h09fa: color = 2'b00;
      13'h09fb: color = 2'b00;
      13'h09fc: color = 2'b11;
      13'h09fd: color = 2'b11;
      13'h09fe: color = 2'b11;
      13'h09ff: color = 2'b11;
      13'h0a00: color = 2'b10;
      13'h0a01: color = 2'b10;
      13'h0a02: color = 2'b11;
      13'h0a03: color = 2'b11;
      13'h0a04: color = 2'b00;
      13'h0a05: color = 2'b00;
      13'h0a06: color = 2'b11;
      13'h0a07: color = 2'b11;
      13'h0a08: color = 2'b11;
      13'h0a09: color = 2'b11;
      13'h0a0a: color = 2'b11;
      13'h0a0b: color = 2'b11;
      13'h0a0c: color = 2'b11;
      13'h0a0d: color = 2'b11;
      13'h0a0e: color = 2'b11;
      13'h0a0f: color = 2'b11;
      13'h0a10: color = 2'b11;
      13'h0a11: color = 2'b11;
      13'h0a12: color = 2'b11;
      13'h0a13: color = 2'b11;
      13'h0a14: color = 2'b11;
      13'h0a15: color = 2'b11;
      13'h0a16: color = 2'b11;
      13'h0a17: color = 2'b11;
      13'h0a18: color = 2'b11;
      13'h0a19: color = 2'b11;
      13'h0a1a: color = 2'b00;
      13'h0a1b: color = 2'b00;
      13'h0a1c: color = 2'b10;
      13'h0a1d: color = 2'b10;
      13'h0a1e: color = 2'b11;
      13'h0a1f: color = 2'b11;
      13'h0a20: color = 2'b00;
      13'h0a21: color = 2'b00;
      13'h0a22: color = 2'b11;
      13'h0a23: color = 2'b11;
      13'h0a24: color = 2'b10;
      13'h0a25: color = 2'b10;
      13'h0a26: color = 2'b10;
      13'h0a27: color = 2'b10;
      13'h0a28: color = 2'b10;
      13'h0a29: color = 2'b10;
      13'h0a2a: color = 2'b10;
      13'h0a2b: color = 2'b10;
      13'h0a2c: color = 2'b10;
      13'h0a2d: color = 2'b10;
      13'h0a2e: color = 2'b10;
      13'h0a2f: color = 2'b10;
      13'h0a30: color = 2'b10;
      13'h0a31: color = 2'b10;
      13'h0a32: color = 2'b10;
      13'h0a33: color = 2'b10;
      13'h0a34: color = 2'b10;
      13'h0a35: color = 2'b10;
      13'h0a36: color = 2'b10;
      13'h0a37: color = 2'b10;
      13'h0a38: color = 2'b10;
      13'h0a39: color = 2'b10;
      13'h0a3a: color = 2'b10;
      13'h0a3b: color = 2'b10;
      13'h0a3c: color = 2'b10;
      13'h0a3d: color = 2'b10;
      13'h0a3e: color = 2'b10;
      13'h0a3f: color = 2'b10;
      13'h0a40: color = 2'b10;
      13'h0a41: color = 2'b10;
      13'h0a42: color = 2'b10;
      13'h0a43: color = 2'b10;
      13'h0a44: color = 2'b10;
      13'h0a45: color = 2'b10;
      13'h0a46: color = 2'b10;
      13'h0a47: color = 2'b10;
      13'h0a48: color = 2'b10;
      13'h0a49: color = 2'b10;
      13'h0a4a: color = 2'b10;
      13'h0a4b: color = 2'b10;
      13'h0a4c: color = 2'b10;
      13'h0a4d: color = 2'b10;
      13'h0a4e: color = 2'b10;
      13'h0a4f: color = 2'b10;
      13'h0a50: color = 2'b10;
      13'h0a51: color = 2'b10;
      13'h0a52: color = 2'b10;
      13'h0a53: color = 2'b10;
      13'h0a54: color = 2'b10;
      13'h0a55: color = 2'b10;
      13'h0a56: color = 2'b10;
      13'h0a57: color = 2'b10;
      13'h0a58: color = 2'b10;
      13'h0a59: color = 2'b10;
      13'h0a5a: color = 2'b10;
      13'h0a5b: color = 2'b10;
      13'h0a5c: color = 2'b01;
      13'h0a5d: color = 2'b01;
      13'h0a5e: color = 2'b00;
      13'h0a5f: color = 2'b00;
      13'h0a60: color = 2'b10;
      13'h0a61: color = 2'b10;
      13'h0a62: color = 2'b11;
      13'h0a63: color = 2'b11;
      13'h0a64: color = 2'b00;
      13'h0a65: color = 2'b00;
      13'h0a66: color = 2'b11;
      13'h0a67: color = 2'b11;
      13'h0a68: color = 2'b11;
      13'h0a69: color = 2'b11;
      13'h0a6a: color = 2'b11;
      13'h0a6b: color = 2'b11;
      13'h0a6c: color = 2'b11;
      13'h0a6d: color = 2'b11;
      13'h0a6e: color = 2'b11;
      13'h0a6f: color = 2'b11;
      13'h0a70: color = 2'b11;
      13'h0a71: color = 2'b11;
      13'h0a72: color = 2'b11;
      13'h0a73: color = 2'b11;
      13'h0a74: color = 2'b11;
      13'h0a75: color = 2'b11;
      13'h0a76: color = 2'b11;
      13'h0a77: color = 2'b11;
      13'h0a78: color = 2'b11;
      13'h0a79: color = 2'b11;
      13'h0a7a: color = 2'b00;
      13'h0a7b: color = 2'b00;
      13'h0a7c: color = 2'b10;
      13'h0a7d: color = 2'b10;
      13'h0a7e: color = 2'b11;
      13'h0a7f: color = 2'b11;
      13'h0a80: color = 2'b10;
      13'h0a81: color = 2'b10;
      13'h0a82: color = 2'b11;
      13'h0a83: color = 2'b11;
      13'h0a84: color = 2'b00;
      13'h0a85: color = 2'b00;
      13'h0a86: color = 2'b11;
      13'h0a87: color = 2'b11;
      13'h0a88: color = 2'b11;
      13'h0a89: color = 2'b11;
      13'h0a8a: color = 2'b11;
      13'h0a8b: color = 2'b11;
      13'h0a8c: color = 2'b11;
      13'h0a8d: color = 2'b11;
      13'h0a8e: color = 2'b11;
      13'h0a8f: color = 2'b11;
      13'h0a90: color = 2'b11;
      13'h0a91: color = 2'b11;
      13'h0a92: color = 2'b11;
      13'h0a93: color = 2'b11;
      13'h0a94: color = 2'b11;
      13'h0a95: color = 2'b11;
      13'h0a96: color = 2'b11;
      13'h0a97: color = 2'b11;
      13'h0a98: color = 2'b11;
      13'h0a99: color = 2'b11;
      13'h0a9a: color = 2'b00;
      13'h0a9b: color = 2'b00;
      13'h0a9c: color = 2'b10;
      13'h0a9d: color = 2'b10;
      13'h0a9e: color = 2'b11;
      13'h0a9f: color = 2'b11;
      13'h0aa0: color = 2'b00;
      13'h0aa1: color = 2'b00;
      13'h0aa2: color = 2'b11;
      13'h0aa3: color = 2'b11;
      13'h0aa4: color = 2'b10;
      13'h0aa5: color = 2'b10;
      13'h0aa6: color = 2'b10;
      13'h0aa7: color = 2'b10;
      13'h0aa8: color = 2'b10;
      13'h0aa9: color = 2'b10;
      13'h0aaa: color = 2'b10;
      13'h0aab: color = 2'b10;
      13'h0aac: color = 2'b10;
      13'h0aad: color = 2'b10;
      13'h0aae: color = 2'b10;
      13'h0aaf: color = 2'b10;
      13'h0ab0: color = 2'b10;
      13'h0ab1: color = 2'b10;
      13'h0ab2: color = 2'b10;
      13'h0ab3: color = 2'b10;
      13'h0ab4: color = 2'b10;
      13'h0ab5: color = 2'b10;
      13'h0ab6: color = 2'b10;
      13'h0ab7: color = 2'b10;
      13'h0ab8: color = 2'b10;
      13'h0ab9: color = 2'b10;
      13'h0aba: color = 2'b10;
      13'h0abb: color = 2'b10;
      13'h0abc: color = 2'b10;
      13'h0abd: color = 2'b10;
      13'h0abe: color = 2'b10;
      13'h0abf: color = 2'b10;
      13'h0ac0: color = 2'b10;
      13'h0ac1: color = 2'b10;
      13'h0ac2: color = 2'b10;
      13'h0ac3: color = 2'b10;
      13'h0ac4: color = 2'b10;
      13'h0ac5: color = 2'b10;
      13'h0ac6: color = 2'b10;
      13'h0ac7: color = 2'b10;
      13'h0ac8: color = 2'b10;
      13'h0ac9: color = 2'b10;
      13'h0aca: color = 2'b10;
      13'h0acb: color = 2'b10;
      13'h0acc: color = 2'b10;
      13'h0acd: color = 2'b10;
      13'h0ace: color = 2'b10;
      13'h0acf: color = 2'b10;
      13'h0ad0: color = 2'b10;
      13'h0ad1: color = 2'b10;
      13'h0ad2: color = 2'b10;
      13'h0ad3: color = 2'b10;
      13'h0ad4: color = 2'b10;
      13'h0ad5: color = 2'b10;
      13'h0ad6: color = 2'b10;
      13'h0ad7: color = 2'b10;
      13'h0ad8: color = 2'b10;
      13'h0ad9: color = 2'b10;
      13'h0ada: color = 2'b10;
      13'h0adb: color = 2'b10;
      13'h0adc: color = 2'b01;
      13'h0add: color = 2'b01;
      13'h0ade: color = 2'b00;
      13'h0adf: color = 2'b00;
      13'h0ae0: color = 2'b10;
      13'h0ae1: color = 2'b10;
      13'h0ae2: color = 2'b11;
      13'h0ae3: color = 2'b11;
      13'h0ae4: color = 2'b00;
      13'h0ae5: color = 2'b00;
      13'h0ae6: color = 2'b11;
      13'h0ae7: color = 2'b11;
      13'h0ae8: color = 2'b11;
      13'h0ae9: color = 2'b11;
      13'h0aea: color = 2'b11;
      13'h0aeb: color = 2'b11;
      13'h0aec: color = 2'b11;
      13'h0aed: color = 2'b11;
      13'h0aee: color = 2'b11;
      13'h0aef: color = 2'b11;
      13'h0af0: color = 2'b11;
      13'h0af1: color = 2'b11;
      13'h0af2: color = 2'b11;
      13'h0af3: color = 2'b11;
      13'h0af4: color = 2'b11;
      13'h0af5: color = 2'b11;
      13'h0af6: color = 2'b11;
      13'h0af7: color = 2'b11;
      13'h0af8: color = 2'b11;
      13'h0af9: color = 2'b11;
      13'h0afa: color = 2'b00;
      13'h0afb: color = 2'b00;
      13'h0afc: color = 2'b10;
      13'h0afd: color = 2'b10;
      13'h0afe: color = 2'b11;
      13'h0aff: color = 2'b11;
      13'h0b00: color = 2'b11;
      13'h0b01: color = 2'b11;
      13'h0b02: color = 2'b11;
      13'h0b03: color = 2'b11;
      13'h0b04: color = 2'b00;
      13'h0b05: color = 2'b00;
      13'h0b06: color = 2'b10;
      13'h0b07: color = 2'b10;
      13'h0b08: color = 2'b10;
      13'h0b09: color = 2'b10;
      13'h0b0a: color = 2'b10;
      13'h0b0b: color = 2'b10;
      13'h0b0c: color = 2'b10;
      13'h0b0d: color = 2'b10;
      13'h0b0e: color = 2'b10;
      13'h0b0f: color = 2'b10;
      13'h0b10: color = 2'b10;
      13'h0b11: color = 2'b10;
      13'h0b12: color = 2'b10;
      13'h0b13: color = 2'b10;
      13'h0b14: color = 2'b10;
      13'h0b15: color = 2'b10;
      13'h0b16: color = 2'b10;
      13'h0b17: color = 2'b10;
      13'h0b18: color = 2'b10;
      13'h0b19: color = 2'b10;
      13'h0b1a: color = 2'b00;
      13'h0b1b: color = 2'b00;
      13'h0b1c: color = 2'b11;
      13'h0b1d: color = 2'b11;
      13'h0b1e: color = 2'b10;
      13'h0b1f: color = 2'b10;
      13'h0b20: color = 2'b00;
      13'h0b21: color = 2'b00;
      13'h0b22: color = 2'b11;
      13'h0b23: color = 2'b11;
      13'h0b24: color = 2'b10;
      13'h0b25: color = 2'b10;
      13'h0b26: color = 2'b10;
      13'h0b27: color = 2'b10;
      13'h0b28: color = 2'b10;
      13'h0b29: color = 2'b10;
      13'h0b2a: color = 2'b10;
      13'h0b2b: color = 2'b10;
      13'h0b2c: color = 2'b10;
      13'h0b2d: color = 2'b10;
      13'h0b2e: color = 2'b10;
      13'h0b2f: color = 2'b10;
      13'h0b30: color = 2'b10;
      13'h0b31: color = 2'b10;
      13'h0b32: color = 2'b10;
      13'h0b33: color = 2'b10;
      13'h0b34: color = 2'b10;
      13'h0b35: color = 2'b10;
      13'h0b36: color = 2'b10;
      13'h0b37: color = 2'b10;
      13'h0b38: color = 2'b10;
      13'h0b39: color = 2'b10;
      13'h0b3a: color = 2'b10;
      13'h0b3b: color = 2'b10;
      13'h0b3c: color = 2'b10;
      13'h0b3d: color = 2'b10;
      13'h0b3e: color = 2'b10;
      13'h0b3f: color = 2'b10;
      13'h0b40: color = 2'b10;
      13'h0b41: color = 2'b10;
      13'h0b42: color = 2'b10;
      13'h0b43: color = 2'b10;
      13'h0b44: color = 2'b10;
      13'h0b45: color = 2'b10;
      13'h0b46: color = 2'b10;
      13'h0b47: color = 2'b10;
      13'h0b48: color = 2'b10;
      13'h0b49: color = 2'b10;
      13'h0b4a: color = 2'b10;
      13'h0b4b: color = 2'b10;
      13'h0b4c: color = 2'b10;
      13'h0b4d: color = 2'b10;
      13'h0b4e: color = 2'b10;
      13'h0b4f: color = 2'b10;
      13'h0b50: color = 2'b10;
      13'h0b51: color = 2'b10;
      13'h0b52: color = 2'b10;
      13'h0b53: color = 2'b10;
      13'h0b54: color = 2'b10;
      13'h0b55: color = 2'b10;
      13'h0b56: color = 2'b10;
      13'h0b57: color = 2'b10;
      13'h0b58: color = 2'b10;
      13'h0b59: color = 2'b10;
      13'h0b5a: color = 2'b10;
      13'h0b5b: color = 2'b10;
      13'h0b5c: color = 2'b01;
      13'h0b5d: color = 2'b01;
      13'h0b5e: color = 2'b00;
      13'h0b5f: color = 2'b00;
      13'h0b60: color = 2'b11;
      13'h0b61: color = 2'b11;
      13'h0b62: color = 2'b11;
      13'h0b63: color = 2'b11;
      13'h0b64: color = 2'b00;
      13'h0b65: color = 2'b00;
      13'h0b66: color = 2'b10;
      13'h0b67: color = 2'b10;
      13'h0b68: color = 2'b10;
      13'h0b69: color = 2'b10;
      13'h0b6a: color = 2'b10;
      13'h0b6b: color = 2'b10;
      13'h0b6c: color = 2'b10;
      13'h0b6d: color = 2'b10;
      13'h0b6e: color = 2'b10;
      13'h0b6f: color = 2'b10;
      13'h0b70: color = 2'b10;
      13'h0b71: color = 2'b10;
      13'h0b72: color = 2'b10;
      13'h0b73: color = 2'b10;
      13'h0b74: color = 2'b10;
      13'h0b75: color = 2'b10;
      13'h0b76: color = 2'b10;
      13'h0b77: color = 2'b10;
      13'h0b78: color = 2'b10;
      13'h0b79: color = 2'b10;
      13'h0b7a: color = 2'b00;
      13'h0b7b: color = 2'b00;
      13'h0b7c: color = 2'b11;
      13'h0b7d: color = 2'b11;
      13'h0b7e: color = 2'b10;
      13'h0b7f: color = 2'b10;
      13'h0b80: color = 2'b11;
      13'h0b81: color = 2'b11;
      13'h0b82: color = 2'b11;
      13'h0b83: color = 2'b11;
      13'h0b84: color = 2'b00;
      13'h0b85: color = 2'b00;
      13'h0b86: color = 2'b10;
      13'h0b87: color = 2'b10;
      13'h0b88: color = 2'b10;
      13'h0b89: color = 2'b10;
      13'h0b8a: color = 2'b10;
      13'h0b8b: color = 2'b10;
      13'h0b8c: color = 2'b10;
      13'h0b8d: color = 2'b10;
      13'h0b8e: color = 2'b10;
      13'h0b8f: color = 2'b10;
      13'h0b90: color = 2'b10;
      13'h0b91: color = 2'b10;
      13'h0b92: color = 2'b10;
      13'h0b93: color = 2'b10;
      13'h0b94: color = 2'b10;
      13'h0b95: color = 2'b10;
      13'h0b96: color = 2'b10;
      13'h0b97: color = 2'b10;
      13'h0b98: color = 2'b10;
      13'h0b99: color = 2'b10;
      13'h0b9a: color = 2'b00;
      13'h0b9b: color = 2'b00;
      13'h0b9c: color = 2'b11;
      13'h0b9d: color = 2'b11;
      13'h0b9e: color = 2'b10;
      13'h0b9f: color = 2'b10;
      13'h0ba0: color = 2'b00;
      13'h0ba1: color = 2'b00;
      13'h0ba2: color = 2'b11;
      13'h0ba3: color = 2'b11;
      13'h0ba4: color = 2'b10;
      13'h0ba5: color = 2'b10;
      13'h0ba6: color = 2'b10;
      13'h0ba7: color = 2'b10;
      13'h0ba8: color = 2'b10;
      13'h0ba9: color = 2'b10;
      13'h0baa: color = 2'b10;
      13'h0bab: color = 2'b10;
      13'h0bac: color = 2'b10;
      13'h0bad: color = 2'b10;
      13'h0bae: color = 2'b10;
      13'h0baf: color = 2'b10;
      13'h0bb0: color = 2'b10;
      13'h0bb1: color = 2'b10;
      13'h0bb2: color = 2'b10;
      13'h0bb3: color = 2'b10;
      13'h0bb4: color = 2'b10;
      13'h0bb5: color = 2'b10;
      13'h0bb6: color = 2'b10;
      13'h0bb7: color = 2'b10;
      13'h0bb8: color = 2'b10;
      13'h0bb9: color = 2'b10;
      13'h0bba: color = 2'b10;
      13'h0bbb: color = 2'b10;
      13'h0bbc: color = 2'b10;
      13'h0bbd: color = 2'b10;
      13'h0bbe: color = 2'b10;
      13'h0bbf: color = 2'b10;
      13'h0bc0: color = 2'b10;
      13'h0bc1: color = 2'b10;
      13'h0bc2: color = 2'b10;
      13'h0bc3: color = 2'b10;
      13'h0bc4: color = 2'b10;
      13'h0bc5: color = 2'b10;
      13'h0bc6: color = 2'b10;
      13'h0bc7: color = 2'b10;
      13'h0bc8: color = 2'b10;
      13'h0bc9: color = 2'b10;
      13'h0bca: color = 2'b10;
      13'h0bcb: color = 2'b10;
      13'h0bcc: color = 2'b10;
      13'h0bcd: color = 2'b10;
      13'h0bce: color = 2'b10;
      13'h0bcf: color = 2'b10;
      13'h0bd0: color = 2'b10;
      13'h0bd1: color = 2'b10;
      13'h0bd2: color = 2'b10;
      13'h0bd3: color = 2'b10;
      13'h0bd4: color = 2'b10;
      13'h0bd5: color = 2'b10;
      13'h0bd6: color = 2'b10;
      13'h0bd7: color = 2'b10;
      13'h0bd8: color = 2'b10;
      13'h0bd9: color = 2'b10;
      13'h0bda: color = 2'b10;
      13'h0bdb: color = 2'b10;
      13'h0bdc: color = 2'b01;
      13'h0bdd: color = 2'b01;
      13'h0bde: color = 2'b00;
      13'h0bdf: color = 2'b00;
      13'h0be0: color = 2'b11;
      13'h0be1: color = 2'b11;
      13'h0be2: color = 2'b11;
      13'h0be3: color = 2'b11;
      13'h0be4: color = 2'b00;
      13'h0be5: color = 2'b00;
      13'h0be6: color = 2'b10;
      13'h0be7: color = 2'b10;
      13'h0be8: color = 2'b10;
      13'h0be9: color = 2'b10;
      13'h0bea: color = 2'b10;
      13'h0beb: color = 2'b10;
      13'h0bec: color = 2'b10;
      13'h0bed: color = 2'b10;
      13'h0bee: color = 2'b10;
      13'h0bef: color = 2'b10;
      13'h0bf0: color = 2'b10;
      13'h0bf1: color = 2'b10;
      13'h0bf2: color = 2'b10;
      13'h0bf3: color = 2'b10;
      13'h0bf4: color = 2'b10;
      13'h0bf5: color = 2'b10;
      13'h0bf6: color = 2'b10;
      13'h0bf7: color = 2'b10;
      13'h0bf8: color = 2'b10;
      13'h0bf9: color = 2'b10;
      13'h0bfa: color = 2'b00;
      13'h0bfb: color = 2'b00;
      13'h0bfc: color = 2'b11;
      13'h0bfd: color = 2'b11;
      13'h0bfe: color = 2'b10;
      13'h0bff: color = 2'b10;
      13'h0c00: color = 2'b10;
      13'h0c01: color = 2'b10;
      13'h0c02: color = 2'b11;
      13'h0c03: color = 2'b11;
      13'h0c04: color = 2'b00;
      13'h0c05: color = 2'b00;
      13'h0c06: color = 2'b10;
      13'h0c07: color = 2'b10;
      13'h0c08: color = 2'b00;
      13'h0c09: color = 2'b00;
      13'h0c0a: color = 2'b00;
      13'h0c0b: color = 2'b00;
      13'h0c0c: color = 2'b00;
      13'h0c0d: color = 2'b00;
      13'h0c0e: color = 2'b00;
      13'h0c0f: color = 2'b00;
      13'h0c10: color = 2'b00;
      13'h0c11: color = 2'b00;
      13'h0c12: color = 2'b00;
      13'h0c13: color = 2'b00;
      13'h0c14: color = 2'b00;
      13'h0c15: color = 2'b00;
      13'h0c16: color = 2'b00;
      13'h0c17: color = 2'b00;
      13'h0c18: color = 2'b10;
      13'h0c19: color = 2'b10;
      13'h0c1a: color = 2'b00;
      13'h0c1b: color = 2'b00;
      13'h0c1c: color = 2'b11;
      13'h0c1d: color = 2'b11;
      13'h0c1e: color = 2'b11;
      13'h0c1f: color = 2'b11;
      13'h0c20: color = 2'b00;
      13'h0c21: color = 2'b00;
      13'h0c22: color = 2'b11;
      13'h0c23: color = 2'b11;
      13'h0c24: color = 2'b10;
      13'h0c25: color = 2'b10;
      13'h0c26: color = 2'b10;
      13'h0c27: color = 2'b10;
      13'h0c28: color = 2'b10;
      13'h0c29: color = 2'b10;
      13'h0c2a: color = 2'b10;
      13'h0c2b: color = 2'b10;
      13'h0c2c: color = 2'b10;
      13'h0c2d: color = 2'b10;
      13'h0c2e: color = 2'b10;
      13'h0c2f: color = 2'b10;
      13'h0c30: color = 2'b10;
      13'h0c31: color = 2'b10;
      13'h0c32: color = 2'b10;
      13'h0c33: color = 2'b10;
      13'h0c34: color = 2'b10;
      13'h0c35: color = 2'b10;
      13'h0c36: color = 2'b10;
      13'h0c37: color = 2'b10;
      13'h0c38: color = 2'b10;
      13'h0c39: color = 2'b10;
      13'h0c3a: color = 2'b10;
      13'h0c3b: color = 2'b10;
      13'h0c3c: color = 2'b10;
      13'h0c3d: color = 2'b10;
      13'h0c3e: color = 2'b10;
      13'h0c3f: color = 2'b10;
      13'h0c40: color = 2'b10;
      13'h0c41: color = 2'b10;
      13'h0c42: color = 2'b10;
      13'h0c43: color = 2'b10;
      13'h0c44: color = 2'b10;
      13'h0c45: color = 2'b10;
      13'h0c46: color = 2'b10;
      13'h0c47: color = 2'b10;
      13'h0c48: color = 2'b10;
      13'h0c49: color = 2'b10;
      13'h0c4a: color = 2'b10;
      13'h0c4b: color = 2'b10;
      13'h0c4c: color = 2'b10;
      13'h0c4d: color = 2'b10;
      13'h0c4e: color = 2'b10;
      13'h0c4f: color = 2'b10;
      13'h0c50: color = 2'b10;
      13'h0c51: color = 2'b10;
      13'h0c52: color = 2'b10;
      13'h0c53: color = 2'b10;
      13'h0c54: color = 2'b10;
      13'h0c55: color = 2'b10;
      13'h0c56: color = 2'b10;
      13'h0c57: color = 2'b10;
      13'h0c58: color = 2'b10;
      13'h0c59: color = 2'b10;
      13'h0c5a: color = 2'b10;
      13'h0c5b: color = 2'b10;
      13'h0c5c: color = 2'b01;
      13'h0c5d: color = 2'b01;
      13'h0c5e: color = 2'b00;
      13'h0c5f: color = 2'b00;
      13'h0c60: color = 2'b10;
      13'h0c61: color = 2'b10;
      13'h0c62: color = 2'b11;
      13'h0c63: color = 2'b11;
      13'h0c64: color = 2'b00;
      13'h0c65: color = 2'b00;
      13'h0c66: color = 2'b10;
      13'h0c67: color = 2'b10;
      13'h0c68: color = 2'b00;
      13'h0c69: color = 2'b00;
      13'h0c6a: color = 2'b00;
      13'h0c6b: color = 2'b00;
      13'h0c6c: color = 2'b00;
      13'h0c6d: color = 2'b00;
      13'h0c6e: color = 2'b00;
      13'h0c6f: color = 2'b00;
      13'h0c70: color = 2'b00;
      13'h0c71: color = 2'b00;
      13'h0c72: color = 2'b00;
      13'h0c73: color = 2'b00;
      13'h0c74: color = 2'b00;
      13'h0c75: color = 2'b00;
      13'h0c76: color = 2'b00;
      13'h0c77: color = 2'b00;
      13'h0c78: color = 2'b10;
      13'h0c79: color = 2'b10;
      13'h0c7a: color = 2'b00;
      13'h0c7b: color = 2'b00;
      13'h0c7c: color = 2'b11;
      13'h0c7d: color = 2'b11;
      13'h0c7e: color = 2'b11;
      13'h0c7f: color = 2'b11;
      13'h0c80: color = 2'b10;
      13'h0c81: color = 2'b10;
      13'h0c82: color = 2'b11;
      13'h0c83: color = 2'b11;
      13'h0c84: color = 2'b00;
      13'h0c85: color = 2'b00;
      13'h0c86: color = 2'b10;
      13'h0c87: color = 2'b10;
      13'h0c88: color = 2'b00;
      13'h0c89: color = 2'b00;
      13'h0c8a: color = 2'b00;
      13'h0c8b: color = 2'b00;
      13'h0c8c: color = 2'b00;
      13'h0c8d: color = 2'b00;
      13'h0c8e: color = 2'b00;
      13'h0c8f: color = 2'b00;
      13'h0c90: color = 2'b00;
      13'h0c91: color = 2'b00;
      13'h0c92: color = 2'b00;
      13'h0c93: color = 2'b00;
      13'h0c94: color = 2'b00;
      13'h0c95: color = 2'b00;
      13'h0c96: color = 2'b00;
      13'h0c97: color = 2'b00;
      13'h0c98: color = 2'b10;
      13'h0c99: color = 2'b10;
      13'h0c9a: color = 2'b00;
      13'h0c9b: color = 2'b00;
      13'h0c9c: color = 2'b11;
      13'h0c9d: color = 2'b11;
      13'h0c9e: color = 2'b11;
      13'h0c9f: color = 2'b11;
      13'h0ca0: color = 2'b00;
      13'h0ca1: color = 2'b00;
      13'h0ca2: color = 2'b11;
      13'h0ca3: color = 2'b11;
      13'h0ca4: color = 2'b10;
      13'h0ca5: color = 2'b10;
      13'h0ca6: color = 2'b10;
      13'h0ca7: color = 2'b10;
      13'h0ca8: color = 2'b10;
      13'h0ca9: color = 2'b10;
      13'h0caa: color = 2'b10;
      13'h0cab: color = 2'b10;
      13'h0cac: color = 2'b10;
      13'h0cad: color = 2'b10;
      13'h0cae: color = 2'b10;
      13'h0caf: color = 2'b10;
      13'h0cb0: color = 2'b10;
      13'h0cb1: color = 2'b10;
      13'h0cb2: color = 2'b10;
      13'h0cb3: color = 2'b10;
      13'h0cb4: color = 2'b10;
      13'h0cb5: color = 2'b10;
      13'h0cb6: color = 2'b10;
      13'h0cb7: color = 2'b10;
      13'h0cb8: color = 2'b10;
      13'h0cb9: color = 2'b10;
      13'h0cba: color = 2'b10;
      13'h0cbb: color = 2'b10;
      13'h0cbc: color = 2'b10;
      13'h0cbd: color = 2'b10;
      13'h0cbe: color = 2'b10;
      13'h0cbf: color = 2'b10;
      13'h0cc0: color = 2'b10;
      13'h0cc1: color = 2'b10;
      13'h0cc2: color = 2'b10;
      13'h0cc3: color = 2'b10;
      13'h0cc4: color = 2'b10;
      13'h0cc5: color = 2'b10;
      13'h0cc6: color = 2'b10;
      13'h0cc7: color = 2'b10;
      13'h0cc8: color = 2'b10;
      13'h0cc9: color = 2'b10;
      13'h0cca: color = 2'b10;
      13'h0ccb: color = 2'b10;
      13'h0ccc: color = 2'b10;
      13'h0ccd: color = 2'b10;
      13'h0cce: color = 2'b10;
      13'h0ccf: color = 2'b10;
      13'h0cd0: color = 2'b10;
      13'h0cd1: color = 2'b10;
      13'h0cd2: color = 2'b10;
      13'h0cd3: color = 2'b10;
      13'h0cd4: color = 2'b10;
      13'h0cd5: color = 2'b10;
      13'h0cd6: color = 2'b10;
      13'h0cd7: color = 2'b10;
      13'h0cd8: color = 2'b10;
      13'h0cd9: color = 2'b10;
      13'h0cda: color = 2'b10;
      13'h0cdb: color = 2'b10;
      13'h0cdc: color = 2'b01;
      13'h0cdd: color = 2'b01;
      13'h0cde: color = 2'b00;
      13'h0cdf: color = 2'b00;
      13'h0ce0: color = 2'b10;
      13'h0ce1: color = 2'b10;
      13'h0ce2: color = 2'b11;
      13'h0ce3: color = 2'b11;
      13'h0ce4: color = 2'b00;
      13'h0ce5: color = 2'b00;
      13'h0ce6: color = 2'b10;
      13'h0ce7: color = 2'b10;
      13'h0ce8: color = 2'b00;
      13'h0ce9: color = 2'b00;
      13'h0cea: color = 2'b00;
      13'h0ceb: color = 2'b00;
      13'h0cec: color = 2'b00;
      13'h0ced: color = 2'b00;
      13'h0cee: color = 2'b00;
      13'h0cef: color = 2'b00;
      13'h0cf0: color = 2'b00;
      13'h0cf1: color = 2'b00;
      13'h0cf2: color = 2'b00;
      13'h0cf3: color = 2'b00;
      13'h0cf4: color = 2'b00;
      13'h0cf5: color = 2'b00;
      13'h0cf6: color = 2'b00;
      13'h0cf7: color = 2'b00;
      13'h0cf8: color = 2'b10;
      13'h0cf9: color = 2'b10;
      13'h0cfa: color = 2'b00;
      13'h0cfb: color = 2'b00;
      13'h0cfc: color = 2'b11;
      13'h0cfd: color = 2'b11;
      13'h0cfe: color = 2'b11;
      13'h0cff: color = 2'b11;
      13'h0d00: color = 2'b11;
      13'h0d01: color = 2'b11;
      13'h0d02: color = 2'b10;
      13'h0d03: color = 2'b10;
      13'h0d04: color = 2'b00;
      13'h0d05: color = 2'b00;
      13'h0d06: color = 2'b10;
      13'h0d07: color = 2'b10;
      13'h0d08: color = 2'b00;
      13'h0d09: color = 2'b00;
      13'h0d0a: color = 2'b11;
      13'h0d0b: color = 2'b11;
      13'h0d0c: color = 2'b11;
      13'h0d0d: color = 2'b11;
      13'h0d0e: color = 2'b11;
      13'h0d0f: color = 2'b11;
      13'h0d10: color = 2'b11;
      13'h0d11: color = 2'b11;
      13'h0d12: color = 2'b10;
      13'h0d13: color = 2'b10;
      13'h0d14: color = 2'b11;
      13'h0d15: color = 2'b11;
      13'h0d16: color = 2'b00;
      13'h0d17: color = 2'b00;
      13'h0d18: color = 2'b10;
      13'h0d19: color = 2'b10;
      13'h0d1a: color = 2'b00;
      13'h0d1b: color = 2'b00;
      13'h0d1c: color = 2'b11;
      13'h0d1d: color = 2'b11;
      13'h0d1e: color = 2'b11;
      13'h0d1f: color = 2'b11;
      13'h0d20: color = 2'b00;
      13'h0d21: color = 2'b00;
      13'h0d22: color = 2'b11;
      13'h0d23: color = 2'b11;
      13'h0d24: color = 2'b10;
      13'h0d25: color = 2'b10;
      13'h0d26: color = 2'b10;
      13'h0d27: color = 2'b10;
      13'h0d28: color = 2'b10;
      13'h0d29: color = 2'b10;
      13'h0d2a: color = 2'b10;
      13'h0d2b: color = 2'b10;
      13'h0d2c: color = 2'b10;
      13'h0d2d: color = 2'b10;
      13'h0d2e: color = 2'b10;
      13'h0d2f: color = 2'b10;
      13'h0d30: color = 2'b10;
      13'h0d31: color = 2'b10;
      13'h0d32: color = 2'b10;
      13'h0d33: color = 2'b10;
      13'h0d34: color = 2'b10;
      13'h0d35: color = 2'b10;
      13'h0d36: color = 2'b10;
      13'h0d37: color = 2'b10;
      13'h0d38: color = 2'b10;
      13'h0d39: color = 2'b10;
      13'h0d3a: color = 2'b10;
      13'h0d3b: color = 2'b10;
      13'h0d3c: color = 2'b10;
      13'h0d3d: color = 2'b10;
      13'h0d3e: color = 2'b10;
      13'h0d3f: color = 2'b10;
      13'h0d40: color = 2'b10;
      13'h0d41: color = 2'b10;
      13'h0d42: color = 2'b10;
      13'h0d43: color = 2'b10;
      13'h0d44: color = 2'b10;
      13'h0d45: color = 2'b10;
      13'h0d46: color = 2'b10;
      13'h0d47: color = 2'b10;
      13'h0d48: color = 2'b10;
      13'h0d49: color = 2'b10;
      13'h0d4a: color = 2'b10;
      13'h0d4b: color = 2'b10;
      13'h0d4c: color = 2'b10;
      13'h0d4d: color = 2'b10;
      13'h0d4e: color = 2'b10;
      13'h0d4f: color = 2'b10;
      13'h0d50: color = 2'b10;
      13'h0d51: color = 2'b10;
      13'h0d52: color = 2'b10;
      13'h0d53: color = 2'b10;
      13'h0d54: color = 2'b10;
      13'h0d55: color = 2'b10;
      13'h0d56: color = 2'b10;
      13'h0d57: color = 2'b10;
      13'h0d58: color = 2'b10;
      13'h0d59: color = 2'b10;
      13'h0d5a: color = 2'b10;
      13'h0d5b: color = 2'b10;
      13'h0d5c: color = 2'b01;
      13'h0d5d: color = 2'b01;
      13'h0d5e: color = 2'b00;
      13'h0d5f: color = 2'b00;
      13'h0d60: color = 2'b11;
      13'h0d61: color = 2'b11;
      13'h0d62: color = 2'b10;
      13'h0d63: color = 2'b10;
      13'h0d64: color = 2'b00;
      13'h0d65: color = 2'b00;
      13'h0d66: color = 2'b10;
      13'h0d67: color = 2'b10;
      13'h0d68: color = 2'b00;
      13'h0d69: color = 2'b00;
      13'h0d6a: color = 2'b11;
      13'h0d6b: color = 2'b11;
      13'h0d6c: color = 2'b11;
      13'h0d6d: color = 2'b11;
      13'h0d6e: color = 2'b11;
      13'h0d6f: color = 2'b11;
      13'h0d70: color = 2'b11;
      13'h0d71: color = 2'b11;
      13'h0d72: color = 2'b10;
      13'h0d73: color = 2'b10;
      13'h0d74: color = 2'b11;
      13'h0d75: color = 2'b11;
      13'h0d76: color = 2'b00;
      13'h0d77: color = 2'b00;
      13'h0d78: color = 2'b10;
      13'h0d79: color = 2'b10;
      13'h0d7a: color = 2'b00;
      13'h0d7b: color = 2'b00;
      13'h0d7c: color = 2'b11;
      13'h0d7d: color = 2'b11;
      13'h0d7e: color = 2'b11;
      13'h0d7f: color = 2'b11;
      13'h0d80: color = 2'b11;
      13'h0d81: color = 2'b11;
      13'h0d82: color = 2'b10;
      13'h0d83: color = 2'b10;
      13'h0d84: color = 2'b00;
      13'h0d85: color = 2'b00;
      13'h0d86: color = 2'b10;
      13'h0d87: color = 2'b10;
      13'h0d88: color = 2'b00;
      13'h0d89: color = 2'b00;
      13'h0d8a: color = 2'b11;
      13'h0d8b: color = 2'b11;
      13'h0d8c: color = 2'b11;
      13'h0d8d: color = 2'b11;
      13'h0d8e: color = 2'b11;
      13'h0d8f: color = 2'b11;
      13'h0d90: color = 2'b11;
      13'h0d91: color = 2'b11;
      13'h0d92: color = 2'b10;
      13'h0d93: color = 2'b10;
      13'h0d94: color = 2'b11;
      13'h0d95: color = 2'b11;
      13'h0d96: color = 2'b00;
      13'h0d97: color = 2'b00;
      13'h0d98: color = 2'b10;
      13'h0d99: color = 2'b10;
      13'h0d9a: color = 2'b00;
      13'h0d9b: color = 2'b00;
      13'h0d9c: color = 2'b11;
      13'h0d9d: color = 2'b11;
      13'h0d9e: color = 2'b11;
      13'h0d9f: color = 2'b11;
      13'h0da0: color = 2'b00;
      13'h0da1: color = 2'b00;
      13'h0da2: color = 2'b11;
      13'h0da3: color = 2'b11;
      13'h0da4: color = 2'b10;
      13'h0da5: color = 2'b10;
      13'h0da6: color = 2'b10;
      13'h0da7: color = 2'b10;
      13'h0da8: color = 2'b10;
      13'h0da9: color = 2'b10;
      13'h0daa: color = 2'b10;
      13'h0dab: color = 2'b10;
      13'h0dac: color = 2'b10;
      13'h0dad: color = 2'b10;
      13'h0dae: color = 2'b10;
      13'h0daf: color = 2'b10;
      13'h0db0: color = 2'b10;
      13'h0db1: color = 2'b10;
      13'h0db2: color = 2'b10;
      13'h0db3: color = 2'b10;
      13'h0db4: color = 2'b10;
      13'h0db5: color = 2'b10;
      13'h0db6: color = 2'b10;
      13'h0db7: color = 2'b10;
      13'h0db8: color = 2'b10;
      13'h0db9: color = 2'b10;
      13'h0dba: color = 2'b10;
      13'h0dbb: color = 2'b10;
      13'h0dbc: color = 2'b10;
      13'h0dbd: color = 2'b10;
      13'h0dbe: color = 2'b10;
      13'h0dbf: color = 2'b10;
      13'h0dc0: color = 2'b10;
      13'h0dc1: color = 2'b10;
      13'h0dc2: color = 2'b10;
      13'h0dc3: color = 2'b10;
      13'h0dc4: color = 2'b10;
      13'h0dc5: color = 2'b10;
      13'h0dc6: color = 2'b10;
      13'h0dc7: color = 2'b10;
      13'h0dc8: color = 2'b10;
      13'h0dc9: color = 2'b10;
      13'h0dca: color = 2'b10;
      13'h0dcb: color = 2'b10;
      13'h0dcc: color = 2'b10;
      13'h0dcd: color = 2'b10;
      13'h0dce: color = 2'b10;
      13'h0dcf: color = 2'b10;
      13'h0dd0: color = 2'b10;
      13'h0dd1: color = 2'b10;
      13'h0dd2: color = 2'b10;
      13'h0dd3: color = 2'b10;
      13'h0dd4: color = 2'b10;
      13'h0dd5: color = 2'b10;
      13'h0dd6: color = 2'b10;
      13'h0dd7: color = 2'b10;
      13'h0dd8: color = 2'b10;
      13'h0dd9: color = 2'b10;
      13'h0dda: color = 2'b10;
      13'h0ddb: color = 2'b10;
      13'h0ddc: color = 2'b01;
      13'h0ddd: color = 2'b01;
      13'h0dde: color = 2'b00;
      13'h0ddf: color = 2'b00;
      13'h0de0: color = 2'b11;
      13'h0de1: color = 2'b11;
      13'h0de2: color = 2'b10;
      13'h0de3: color = 2'b10;
      13'h0de4: color = 2'b00;
      13'h0de5: color = 2'b00;
      13'h0de6: color = 2'b10;
      13'h0de7: color = 2'b10;
      13'h0de8: color = 2'b00;
      13'h0de9: color = 2'b00;
      13'h0dea: color = 2'b11;
      13'h0deb: color = 2'b11;
      13'h0dec: color = 2'b11;
      13'h0ded: color = 2'b11;
      13'h0dee: color = 2'b11;
      13'h0def: color = 2'b11;
      13'h0df0: color = 2'b11;
      13'h0df1: color = 2'b11;
      13'h0df2: color = 2'b10;
      13'h0df3: color = 2'b10;
      13'h0df4: color = 2'b11;
      13'h0df5: color = 2'b11;
      13'h0df6: color = 2'b00;
      13'h0df7: color = 2'b00;
      13'h0df8: color = 2'b10;
      13'h0df9: color = 2'b10;
      13'h0dfa: color = 2'b00;
      13'h0dfb: color = 2'b00;
      13'h0dfc: color = 2'b11;
      13'h0dfd: color = 2'b11;
      13'h0dfe: color = 2'b11;
      13'h0dff: color = 2'b11;
      13'h0e00: color = 2'b11;
      13'h0e01: color = 2'b11;
      13'h0e02: color = 2'b11;
      13'h0e03: color = 2'b11;
      13'h0e04: color = 2'b00;
      13'h0e05: color = 2'b00;
      13'h0e06: color = 2'b10;
      13'h0e07: color = 2'b10;
      13'h0e08: color = 2'b00;
      13'h0e09: color = 2'b00;
      13'h0e0a: color = 2'b11;
      13'h0e0b: color = 2'b11;
      13'h0e0c: color = 2'b11;
      13'h0e0d: color = 2'b11;
      13'h0e0e: color = 2'b11;
      13'h0e0f: color = 2'b11;
      13'h0e10: color = 2'b11;
      13'h0e11: color = 2'b11;
      13'h0e12: color = 2'b11;
      13'h0e13: color = 2'b11;
      13'h0e14: color = 2'b10;
      13'h0e15: color = 2'b10;
      13'h0e16: color = 2'b00;
      13'h0e17: color = 2'b00;
      13'h0e18: color = 2'b10;
      13'h0e19: color = 2'b10;
      13'h0e1a: color = 2'b00;
      13'h0e1b: color = 2'b00;
      13'h0e1c: color = 2'b11;
      13'h0e1d: color = 2'b11;
      13'h0e1e: color = 2'b11;
      13'h0e1f: color = 2'b11;
      13'h0e20: color = 2'b00;
      13'h0e21: color = 2'b00;
      13'h0e22: color = 2'b11;
      13'h0e23: color = 2'b11;
      13'h0e24: color = 2'b10;
      13'h0e25: color = 2'b10;
      13'h0e26: color = 2'b10;
      13'h0e27: color = 2'b10;
      13'h0e28: color = 2'b10;
      13'h0e29: color = 2'b10;
      13'h0e2a: color = 2'b10;
      13'h0e2b: color = 2'b10;
      13'h0e2c: color = 2'b10;
      13'h0e2d: color = 2'b10;
      13'h0e2e: color = 2'b10;
      13'h0e2f: color = 2'b10;
      13'h0e30: color = 2'b10;
      13'h0e31: color = 2'b10;
      13'h0e32: color = 2'b10;
      13'h0e33: color = 2'b10;
      13'h0e34: color = 2'b10;
      13'h0e35: color = 2'b10;
      13'h0e36: color = 2'b10;
      13'h0e37: color = 2'b10;
      13'h0e38: color = 2'b10;
      13'h0e39: color = 2'b10;
      13'h0e3a: color = 2'b10;
      13'h0e3b: color = 2'b10;
      13'h0e3c: color = 2'b10;
      13'h0e3d: color = 2'b10;
      13'h0e3e: color = 2'b10;
      13'h0e3f: color = 2'b10;
      13'h0e40: color = 2'b10;
      13'h0e41: color = 2'b10;
      13'h0e42: color = 2'b10;
      13'h0e43: color = 2'b10;
      13'h0e44: color = 2'b10;
      13'h0e45: color = 2'b10;
      13'h0e46: color = 2'b10;
      13'h0e47: color = 2'b10;
      13'h0e48: color = 2'b10;
      13'h0e49: color = 2'b10;
      13'h0e4a: color = 2'b10;
      13'h0e4b: color = 2'b10;
      13'h0e4c: color = 2'b10;
      13'h0e4d: color = 2'b10;
      13'h0e4e: color = 2'b10;
      13'h0e4f: color = 2'b10;
      13'h0e50: color = 2'b10;
      13'h0e51: color = 2'b10;
      13'h0e52: color = 2'b10;
      13'h0e53: color = 2'b10;
      13'h0e54: color = 2'b10;
      13'h0e55: color = 2'b10;
      13'h0e56: color = 2'b10;
      13'h0e57: color = 2'b10;
      13'h0e58: color = 2'b10;
      13'h0e59: color = 2'b10;
      13'h0e5a: color = 2'b10;
      13'h0e5b: color = 2'b10;
      13'h0e5c: color = 2'b01;
      13'h0e5d: color = 2'b01;
      13'h0e5e: color = 2'b00;
      13'h0e5f: color = 2'b00;
      13'h0e60: color = 2'b11;
      13'h0e61: color = 2'b11;
      13'h0e62: color = 2'b11;
      13'h0e63: color = 2'b11;
      13'h0e64: color = 2'b00;
      13'h0e65: color = 2'b00;
      13'h0e66: color = 2'b10;
      13'h0e67: color = 2'b10;
      13'h0e68: color = 2'b00;
      13'h0e69: color = 2'b00;
      13'h0e6a: color = 2'b11;
      13'h0e6b: color = 2'b11;
      13'h0e6c: color = 2'b11;
      13'h0e6d: color = 2'b11;
      13'h0e6e: color = 2'b11;
      13'h0e6f: color = 2'b11;
      13'h0e70: color = 2'b11;
      13'h0e71: color = 2'b11;
      13'h0e72: color = 2'b11;
      13'h0e73: color = 2'b11;
      13'h0e74: color = 2'b10;
      13'h0e75: color = 2'b10;
      13'h0e76: color = 2'b00;
      13'h0e77: color = 2'b00;
      13'h0e78: color = 2'b10;
      13'h0e79: color = 2'b10;
      13'h0e7a: color = 2'b00;
      13'h0e7b: color = 2'b00;
      13'h0e7c: color = 2'b11;
      13'h0e7d: color = 2'b11;
      13'h0e7e: color = 2'b11;
      13'h0e7f: color = 2'b11;
      13'h0e80: color = 2'b11;
      13'h0e81: color = 2'b11;
      13'h0e82: color = 2'b11;
      13'h0e83: color = 2'b11;
      13'h0e84: color = 2'b00;
      13'h0e85: color = 2'b00;
      13'h0e86: color = 2'b10;
      13'h0e87: color = 2'b10;
      13'h0e88: color = 2'b00;
      13'h0e89: color = 2'b00;
      13'h0e8a: color = 2'b11;
      13'h0e8b: color = 2'b11;
      13'h0e8c: color = 2'b11;
      13'h0e8d: color = 2'b11;
      13'h0e8e: color = 2'b11;
      13'h0e8f: color = 2'b11;
      13'h0e90: color = 2'b11;
      13'h0e91: color = 2'b11;
      13'h0e92: color = 2'b11;
      13'h0e93: color = 2'b11;
      13'h0e94: color = 2'b10;
      13'h0e95: color = 2'b10;
      13'h0e96: color = 2'b00;
      13'h0e97: color = 2'b00;
      13'h0e98: color = 2'b10;
      13'h0e99: color = 2'b10;
      13'h0e9a: color = 2'b00;
      13'h0e9b: color = 2'b00;
      13'h0e9c: color = 2'b11;
      13'h0e9d: color = 2'b11;
      13'h0e9e: color = 2'b11;
      13'h0e9f: color = 2'b11;
      13'h0ea0: color = 2'b00;
      13'h0ea1: color = 2'b00;
      13'h0ea2: color = 2'b11;
      13'h0ea3: color = 2'b11;
      13'h0ea4: color = 2'b10;
      13'h0ea5: color = 2'b10;
      13'h0ea6: color = 2'b10;
      13'h0ea7: color = 2'b10;
      13'h0ea8: color = 2'b10;
      13'h0ea9: color = 2'b10;
      13'h0eaa: color = 2'b10;
      13'h0eab: color = 2'b10;
      13'h0eac: color = 2'b10;
      13'h0ead: color = 2'b10;
      13'h0eae: color = 2'b10;
      13'h0eaf: color = 2'b10;
      13'h0eb0: color = 2'b10;
      13'h0eb1: color = 2'b10;
      13'h0eb2: color = 2'b10;
      13'h0eb3: color = 2'b10;
      13'h0eb4: color = 2'b10;
      13'h0eb5: color = 2'b10;
      13'h0eb6: color = 2'b10;
      13'h0eb7: color = 2'b10;
      13'h0eb8: color = 2'b10;
      13'h0eb9: color = 2'b10;
      13'h0eba: color = 2'b10;
      13'h0ebb: color = 2'b10;
      13'h0ebc: color = 2'b10;
      13'h0ebd: color = 2'b10;
      13'h0ebe: color = 2'b10;
      13'h0ebf: color = 2'b10;
      13'h0ec0: color = 2'b10;
      13'h0ec1: color = 2'b10;
      13'h0ec2: color = 2'b10;
      13'h0ec3: color = 2'b10;
      13'h0ec4: color = 2'b10;
      13'h0ec5: color = 2'b10;
      13'h0ec6: color = 2'b10;
      13'h0ec7: color = 2'b10;
      13'h0ec8: color = 2'b10;
      13'h0ec9: color = 2'b10;
      13'h0eca: color = 2'b10;
      13'h0ecb: color = 2'b10;
      13'h0ecc: color = 2'b10;
      13'h0ecd: color = 2'b10;
      13'h0ece: color = 2'b10;
      13'h0ecf: color = 2'b10;
      13'h0ed0: color = 2'b10;
      13'h0ed1: color = 2'b10;
      13'h0ed2: color = 2'b10;
      13'h0ed3: color = 2'b10;
      13'h0ed4: color = 2'b10;
      13'h0ed5: color = 2'b10;
      13'h0ed6: color = 2'b10;
      13'h0ed7: color = 2'b10;
      13'h0ed8: color = 2'b10;
      13'h0ed9: color = 2'b10;
      13'h0eda: color = 2'b10;
      13'h0edb: color = 2'b10;
      13'h0edc: color = 2'b01;
      13'h0edd: color = 2'b01;
      13'h0ede: color = 2'b00;
      13'h0edf: color = 2'b00;
      13'h0ee0: color = 2'b11;
      13'h0ee1: color = 2'b11;
      13'h0ee2: color = 2'b11;
      13'h0ee3: color = 2'b11;
      13'h0ee4: color = 2'b00;
      13'h0ee5: color = 2'b00;
      13'h0ee6: color = 2'b10;
      13'h0ee7: color = 2'b10;
      13'h0ee8: color = 2'b00;
      13'h0ee9: color = 2'b00;
      13'h0eea: color = 2'b11;
      13'h0eeb: color = 2'b11;
      13'h0eec: color = 2'b11;
      13'h0eed: color = 2'b11;
      13'h0eee: color = 2'b11;
      13'h0eef: color = 2'b11;
      13'h0ef0: color = 2'b11;
      13'h0ef1: color = 2'b11;
      13'h0ef2: color = 2'b11;
      13'h0ef3: color = 2'b11;
      13'h0ef4: color = 2'b10;
      13'h0ef5: color = 2'b10;
      13'h0ef6: color = 2'b00;
      13'h0ef7: color = 2'b00;
      13'h0ef8: color = 2'b10;
      13'h0ef9: color = 2'b10;
      13'h0efa: color = 2'b00;
      13'h0efb: color = 2'b00;
      13'h0efc: color = 2'b11;
      13'h0efd: color = 2'b11;
      13'h0efe: color = 2'b11;
      13'h0eff: color = 2'b11;
      13'h0f00: color = 2'b11;
      13'h0f01: color = 2'b11;
      13'h0f02: color = 2'b11;
      13'h0f03: color = 2'b11;
      13'h0f04: color = 2'b00;
      13'h0f05: color = 2'b00;
      13'h0f06: color = 2'b00;
      13'h0f07: color = 2'b00;
      13'h0f08: color = 2'b00;
      13'h0f09: color = 2'b00;
      13'h0f0a: color = 2'b11;
      13'h0f0b: color = 2'b11;
      13'h0f0c: color = 2'b11;
      13'h0f0d: color = 2'b11;
      13'h0f0e: color = 2'b11;
      13'h0f0f: color = 2'b11;
      13'h0f10: color = 2'b11;
      13'h0f11: color = 2'b11;
      13'h0f12: color = 2'b11;
      13'h0f13: color = 2'b11;
      13'h0f14: color = 2'b11;
      13'h0f15: color = 2'b11;
      13'h0f16: color = 2'b00;
      13'h0f17: color = 2'b00;
      13'h0f18: color = 2'b00;
      13'h0f19: color = 2'b00;
      13'h0f1a: color = 2'b00;
      13'h0f1b: color = 2'b00;
      13'h0f1c: color = 2'b11;
      13'h0f1d: color = 2'b11;
      13'h0f1e: color = 2'b11;
      13'h0f1f: color = 2'b11;
      13'h0f20: color = 2'b00;
      13'h0f21: color = 2'b00;
      13'h0f22: color = 2'b11;
      13'h0f23: color = 2'b11;
      13'h0f24: color = 2'b10;
      13'h0f25: color = 2'b10;
      13'h0f26: color = 2'b10;
      13'h0f27: color = 2'b10;
      13'h0f28: color = 2'b10;
      13'h0f29: color = 2'b10;
      13'h0f2a: color = 2'b10;
      13'h0f2b: color = 2'b10;
      13'h0f2c: color = 2'b10;
      13'h0f2d: color = 2'b10;
      13'h0f2e: color = 2'b10;
      13'h0f2f: color = 2'b10;
      13'h0f30: color = 2'b10;
      13'h0f31: color = 2'b10;
      13'h0f32: color = 2'b10;
      13'h0f33: color = 2'b10;
      13'h0f34: color = 2'b10;
      13'h0f35: color = 2'b10;
      13'h0f36: color = 2'b10;
      13'h0f37: color = 2'b10;
      13'h0f38: color = 2'b10;
      13'h0f39: color = 2'b10;
      13'h0f3a: color = 2'b10;
      13'h0f3b: color = 2'b10;
      13'h0f3c: color = 2'b10;
      13'h0f3d: color = 2'b10;
      13'h0f3e: color = 2'b10;
      13'h0f3f: color = 2'b10;
      13'h0f40: color = 2'b10;
      13'h0f41: color = 2'b10;
      13'h0f42: color = 2'b10;
      13'h0f43: color = 2'b10;
      13'h0f44: color = 2'b10;
      13'h0f45: color = 2'b10;
      13'h0f46: color = 2'b10;
      13'h0f47: color = 2'b10;
      13'h0f48: color = 2'b10;
      13'h0f49: color = 2'b10;
      13'h0f4a: color = 2'b10;
      13'h0f4b: color = 2'b10;
      13'h0f4c: color = 2'b10;
      13'h0f4d: color = 2'b10;
      13'h0f4e: color = 2'b10;
      13'h0f4f: color = 2'b10;
      13'h0f50: color = 2'b10;
      13'h0f51: color = 2'b10;
      13'h0f52: color = 2'b10;
      13'h0f53: color = 2'b10;
      13'h0f54: color = 2'b10;
      13'h0f55: color = 2'b10;
      13'h0f56: color = 2'b10;
      13'h0f57: color = 2'b10;
      13'h0f58: color = 2'b10;
      13'h0f59: color = 2'b10;
      13'h0f5a: color = 2'b10;
      13'h0f5b: color = 2'b10;
      13'h0f5c: color = 2'b01;
      13'h0f5d: color = 2'b01;
      13'h0f5e: color = 2'b00;
      13'h0f5f: color = 2'b00;
      13'h0f60: color = 2'b11;
      13'h0f61: color = 2'b11;
      13'h0f62: color = 2'b11;
      13'h0f63: color = 2'b11;
      13'h0f64: color = 2'b00;
      13'h0f65: color = 2'b00;
      13'h0f66: color = 2'b00;
      13'h0f67: color = 2'b00;
      13'h0f68: color = 2'b00;
      13'h0f69: color = 2'b00;
      13'h0f6a: color = 2'b11;
      13'h0f6b: color = 2'b11;
      13'h0f6c: color = 2'b11;
      13'h0f6d: color = 2'b11;
      13'h0f6e: color = 2'b11;
      13'h0f6f: color = 2'b11;
      13'h0f70: color = 2'b11;
      13'h0f71: color = 2'b11;
      13'h0f72: color = 2'b11;
      13'h0f73: color = 2'b11;
      13'h0f74: color = 2'b11;
      13'h0f75: color = 2'b11;
      13'h0f76: color = 2'b00;
      13'h0f77: color = 2'b00;
      13'h0f78: color = 2'b00;
      13'h0f79: color = 2'b00;
      13'h0f7a: color = 2'b00;
      13'h0f7b: color = 2'b00;
      13'h0f7c: color = 2'b11;
      13'h0f7d: color = 2'b11;
      13'h0f7e: color = 2'b11;
      13'h0f7f: color = 2'b11;
      13'h0f80: color = 2'b11;
      13'h0f81: color = 2'b11;
      13'h0f82: color = 2'b11;
      13'h0f83: color = 2'b11;
      13'h0f84: color = 2'b00;
      13'h0f85: color = 2'b00;
      13'h0f86: color = 2'b00;
      13'h0f87: color = 2'b00;
      13'h0f88: color = 2'b00;
      13'h0f89: color = 2'b00;
      13'h0f8a: color = 2'b11;
      13'h0f8b: color = 2'b11;
      13'h0f8c: color = 2'b11;
      13'h0f8d: color = 2'b11;
      13'h0f8e: color = 2'b11;
      13'h0f8f: color = 2'b11;
      13'h0f90: color = 2'b11;
      13'h0f91: color = 2'b11;
      13'h0f92: color = 2'b11;
      13'h0f93: color = 2'b11;
      13'h0f94: color = 2'b11;
      13'h0f95: color = 2'b11;
      13'h0f96: color = 2'b00;
      13'h0f97: color = 2'b00;
      13'h0f98: color = 2'b00;
      13'h0f99: color = 2'b00;
      13'h0f9a: color = 2'b00;
      13'h0f9b: color = 2'b00;
      13'h0f9c: color = 2'b11;
      13'h0f9d: color = 2'b11;
      13'h0f9e: color = 2'b11;
      13'h0f9f: color = 2'b11;
      13'h0fa0: color = 2'b00;
      13'h0fa1: color = 2'b00;
      13'h0fa2: color = 2'b11;
      13'h0fa3: color = 2'b11;
      13'h0fa4: color = 2'b10;
      13'h0fa5: color = 2'b10;
      13'h0fa6: color = 2'b10;
      13'h0fa7: color = 2'b10;
      13'h0fa8: color = 2'b10;
      13'h0fa9: color = 2'b10;
      13'h0faa: color = 2'b10;
      13'h0fab: color = 2'b10;
      13'h0fac: color = 2'b10;
      13'h0fad: color = 2'b10;
      13'h0fae: color = 2'b10;
      13'h0faf: color = 2'b10;
      13'h0fb0: color = 2'b10;
      13'h0fb1: color = 2'b10;
      13'h0fb2: color = 2'b10;
      13'h0fb3: color = 2'b10;
      13'h0fb4: color = 2'b10;
      13'h0fb5: color = 2'b10;
      13'h0fb6: color = 2'b10;
      13'h0fb7: color = 2'b10;
      13'h0fb8: color = 2'b10;
      13'h0fb9: color = 2'b10;
      13'h0fba: color = 2'b10;
      13'h0fbb: color = 2'b10;
      13'h0fbc: color = 2'b10;
      13'h0fbd: color = 2'b10;
      13'h0fbe: color = 2'b10;
      13'h0fbf: color = 2'b10;
      13'h0fc0: color = 2'b10;
      13'h0fc1: color = 2'b10;
      13'h0fc2: color = 2'b10;
      13'h0fc3: color = 2'b10;
      13'h0fc4: color = 2'b10;
      13'h0fc5: color = 2'b10;
      13'h0fc6: color = 2'b10;
      13'h0fc7: color = 2'b10;
      13'h0fc8: color = 2'b10;
      13'h0fc9: color = 2'b10;
      13'h0fca: color = 2'b10;
      13'h0fcb: color = 2'b10;
      13'h0fcc: color = 2'b10;
      13'h0fcd: color = 2'b10;
      13'h0fce: color = 2'b10;
      13'h0fcf: color = 2'b10;
      13'h0fd0: color = 2'b10;
      13'h0fd1: color = 2'b10;
      13'h0fd2: color = 2'b10;
      13'h0fd3: color = 2'b10;
      13'h0fd4: color = 2'b10;
      13'h0fd5: color = 2'b10;
      13'h0fd6: color = 2'b10;
      13'h0fd7: color = 2'b10;
      13'h0fd8: color = 2'b10;
      13'h0fd9: color = 2'b10;
      13'h0fda: color = 2'b10;
      13'h0fdb: color = 2'b10;
      13'h0fdc: color = 2'b01;
      13'h0fdd: color = 2'b01;
      13'h0fde: color = 2'b00;
      13'h0fdf: color = 2'b00;
      13'h0fe0: color = 2'b11;
      13'h0fe1: color = 2'b11;
      13'h0fe2: color = 2'b11;
      13'h0fe3: color = 2'b11;
      13'h0fe4: color = 2'b00;
      13'h0fe5: color = 2'b00;
      13'h0fe6: color = 2'b00;
      13'h0fe7: color = 2'b00;
      13'h0fe8: color = 2'b00;
      13'h0fe9: color = 2'b00;
      13'h0fea: color = 2'b11;
      13'h0feb: color = 2'b11;
      13'h0fec: color = 2'b11;
      13'h0fed: color = 2'b11;
      13'h0fee: color = 2'b11;
      13'h0fef: color = 2'b11;
      13'h0ff0: color = 2'b11;
      13'h0ff1: color = 2'b11;
      13'h0ff2: color = 2'b11;
      13'h0ff3: color = 2'b11;
      13'h0ff4: color = 2'b11;
      13'h0ff5: color = 2'b11;
      13'h0ff6: color = 2'b00;
      13'h0ff7: color = 2'b00;
      13'h0ff8: color = 2'b00;
      13'h0ff9: color = 2'b00;
      13'h0ffa: color = 2'b00;
      13'h0ffb: color = 2'b00;
      13'h0ffc: color = 2'b11;
      13'h0ffd: color = 2'b11;
      13'h0ffe: color = 2'b11;
      13'h0fff: color = 2'b11;
      13'h1000: color = 2'b11;
      13'h1001: color = 2'b11;
      13'h1002: color = 2'b11;
      13'h1003: color = 2'b11;
      13'h1004: color = 2'b10;
      13'h1005: color = 2'b10;
      13'h1006: color = 2'b11;
      13'h1007: color = 2'b11;
      13'h1008: color = 2'b10;
      13'h1009: color = 2'b10;
      13'h100a: color = 2'b11;
      13'h100b: color = 2'b11;
      13'h100c: color = 2'b11;
      13'h100d: color = 2'b11;
      13'h100e: color = 2'b11;
      13'h100f: color = 2'b11;
      13'h1010: color = 2'b11;
      13'h1011: color = 2'b11;
      13'h1012: color = 2'b11;
      13'h1013: color = 2'b11;
      13'h1014: color = 2'b10;
      13'h1015: color = 2'b10;
      13'h1016: color = 2'b11;
      13'h1017: color = 2'b11;
      13'h1018: color = 2'b10;
      13'h1019: color = 2'b10;
      13'h101a: color = 2'b11;
      13'h101b: color = 2'b11;
      13'h101c: color = 2'b11;
      13'h101d: color = 2'b11;
      13'h101e: color = 2'b11;
      13'h101f: color = 2'b11;
      13'h1020: color = 2'b00;
      13'h1021: color = 2'b00;
      13'h1022: color = 2'b11;
      13'h1023: color = 2'b11;
      13'h1024: color = 2'b10;
      13'h1025: color = 2'b10;
      13'h1026: color = 2'b10;
      13'h1027: color = 2'b10;
      13'h1028: color = 2'b10;
      13'h1029: color = 2'b10;
      13'h102a: color = 2'b10;
      13'h102b: color = 2'b10;
      13'h102c: color = 2'b10;
      13'h102d: color = 2'b10;
      13'h102e: color = 2'b10;
      13'h102f: color = 2'b10;
      13'h1030: color = 2'b10;
      13'h1031: color = 2'b10;
      13'h1032: color = 2'b10;
      13'h1033: color = 2'b10;
      13'h1034: color = 2'b10;
      13'h1035: color = 2'b10;
      13'h1036: color = 2'b10;
      13'h1037: color = 2'b10;
      13'h1038: color = 2'b10;
      13'h1039: color = 2'b10;
      13'h103a: color = 2'b10;
      13'h103b: color = 2'b10;
      13'h103c: color = 2'b10;
      13'h103d: color = 2'b10;
      13'h103e: color = 2'b10;
      13'h103f: color = 2'b10;
      13'h1040: color = 2'b10;
      13'h1041: color = 2'b10;
      13'h1042: color = 2'b10;
      13'h1043: color = 2'b10;
      13'h1044: color = 2'b10;
      13'h1045: color = 2'b10;
      13'h1046: color = 2'b10;
      13'h1047: color = 2'b10;
      13'h1048: color = 2'b10;
      13'h1049: color = 2'b10;
      13'h104a: color = 2'b10;
      13'h104b: color = 2'b10;
      13'h104c: color = 2'b10;
      13'h104d: color = 2'b10;
      13'h104e: color = 2'b10;
      13'h104f: color = 2'b10;
      13'h1050: color = 2'b10;
      13'h1051: color = 2'b10;
      13'h1052: color = 2'b10;
      13'h1053: color = 2'b10;
      13'h1054: color = 2'b10;
      13'h1055: color = 2'b10;
      13'h1056: color = 2'b10;
      13'h1057: color = 2'b10;
      13'h1058: color = 2'b10;
      13'h1059: color = 2'b10;
      13'h105a: color = 2'b10;
      13'h105b: color = 2'b10;
      13'h105c: color = 2'b01;
      13'h105d: color = 2'b01;
      13'h105e: color = 2'b00;
      13'h105f: color = 2'b00;
      13'h1060: color = 2'b11;
      13'h1061: color = 2'b11;
      13'h1062: color = 2'b11;
      13'h1063: color = 2'b11;
      13'h1064: color = 2'b10;
      13'h1065: color = 2'b10;
      13'h1066: color = 2'b11;
      13'h1067: color = 2'b11;
      13'h1068: color = 2'b10;
      13'h1069: color = 2'b10;
      13'h106a: color = 2'b11;
      13'h106b: color = 2'b11;
      13'h106c: color = 2'b11;
      13'h106d: color = 2'b11;
      13'h106e: color = 2'b11;
      13'h106f: color = 2'b11;
      13'h1070: color = 2'b11;
      13'h1071: color = 2'b11;
      13'h1072: color = 2'b11;
      13'h1073: color = 2'b11;
      13'h1074: color = 2'b10;
      13'h1075: color = 2'b10;
      13'h1076: color = 2'b11;
      13'h1077: color = 2'b11;
      13'h1078: color = 2'b10;
      13'h1079: color = 2'b10;
      13'h107a: color = 2'b11;
      13'h107b: color = 2'b11;
      13'h107c: color = 2'b11;
      13'h107d: color = 2'b11;
      13'h107e: color = 2'b11;
      13'h107f: color = 2'b11;
      13'h1080: color = 2'b11;
      13'h1081: color = 2'b11;
      13'h1082: color = 2'b11;
      13'h1083: color = 2'b11;
      13'h1084: color = 2'b10;
      13'h1085: color = 2'b10;
      13'h1086: color = 2'b11;
      13'h1087: color = 2'b11;
      13'h1088: color = 2'b10;
      13'h1089: color = 2'b10;
      13'h108a: color = 2'b11;
      13'h108b: color = 2'b11;
      13'h108c: color = 2'b11;
      13'h108d: color = 2'b11;
      13'h108e: color = 2'b11;
      13'h108f: color = 2'b11;
      13'h1090: color = 2'b11;
      13'h1091: color = 2'b11;
      13'h1092: color = 2'b11;
      13'h1093: color = 2'b11;
      13'h1094: color = 2'b10;
      13'h1095: color = 2'b10;
      13'h1096: color = 2'b11;
      13'h1097: color = 2'b11;
      13'h1098: color = 2'b10;
      13'h1099: color = 2'b10;
      13'h109a: color = 2'b11;
      13'h109b: color = 2'b11;
      13'h109c: color = 2'b11;
      13'h109d: color = 2'b11;
      13'h109e: color = 2'b11;
      13'h109f: color = 2'b11;
      13'h10a0: color = 2'b00;
      13'h10a1: color = 2'b00;
      13'h10a2: color = 2'b11;
      13'h10a3: color = 2'b11;
      13'h10a4: color = 2'b10;
      13'h10a5: color = 2'b10;
      13'h10a6: color = 2'b10;
      13'h10a7: color = 2'b10;
      13'h10a8: color = 2'b10;
      13'h10a9: color = 2'b10;
      13'h10aa: color = 2'b10;
      13'h10ab: color = 2'b10;
      13'h10ac: color = 2'b10;
      13'h10ad: color = 2'b10;
      13'h10ae: color = 2'b10;
      13'h10af: color = 2'b10;
      13'h10b0: color = 2'b10;
      13'h10b1: color = 2'b10;
      13'h10b2: color = 2'b10;
      13'h10b3: color = 2'b10;
      13'h10b4: color = 2'b10;
      13'h10b5: color = 2'b10;
      13'h10b6: color = 2'b10;
      13'h10b7: color = 2'b10;
      13'h10b8: color = 2'b10;
      13'h10b9: color = 2'b10;
      13'h10ba: color = 2'b10;
      13'h10bb: color = 2'b10;
      13'h10bc: color = 2'b10;
      13'h10bd: color = 2'b10;
      13'h10be: color = 2'b10;
      13'h10bf: color = 2'b10;
      13'h10c0: color = 2'b10;
      13'h10c1: color = 2'b10;
      13'h10c2: color = 2'b10;
      13'h10c3: color = 2'b10;
      13'h10c4: color = 2'b10;
      13'h10c5: color = 2'b10;
      13'h10c6: color = 2'b10;
      13'h10c7: color = 2'b10;
      13'h10c8: color = 2'b10;
      13'h10c9: color = 2'b10;
      13'h10ca: color = 2'b10;
      13'h10cb: color = 2'b10;
      13'h10cc: color = 2'b10;
      13'h10cd: color = 2'b10;
      13'h10ce: color = 2'b10;
      13'h10cf: color = 2'b10;
      13'h10d0: color = 2'b10;
      13'h10d1: color = 2'b10;
      13'h10d2: color = 2'b10;
      13'h10d3: color = 2'b10;
      13'h10d4: color = 2'b10;
      13'h10d5: color = 2'b10;
      13'h10d6: color = 2'b10;
      13'h10d7: color = 2'b10;
      13'h10d8: color = 2'b10;
      13'h10d9: color = 2'b10;
      13'h10da: color = 2'b10;
      13'h10db: color = 2'b10;
      13'h10dc: color = 2'b01;
      13'h10dd: color = 2'b01;
      13'h10de: color = 2'b00;
      13'h10df: color = 2'b00;
      13'h10e0: color = 2'b11;
      13'h10e1: color = 2'b11;
      13'h10e2: color = 2'b11;
      13'h10e3: color = 2'b11;
      13'h10e4: color = 2'b10;
      13'h10e5: color = 2'b10;
      13'h10e6: color = 2'b11;
      13'h10e7: color = 2'b11;
      13'h10e8: color = 2'b10;
      13'h10e9: color = 2'b10;
      13'h10ea: color = 2'b11;
      13'h10eb: color = 2'b11;
      13'h10ec: color = 2'b11;
      13'h10ed: color = 2'b11;
      13'h10ee: color = 2'b11;
      13'h10ef: color = 2'b11;
      13'h10f0: color = 2'b11;
      13'h10f1: color = 2'b11;
      13'h10f2: color = 2'b11;
      13'h10f3: color = 2'b11;
      13'h10f4: color = 2'b10;
      13'h10f5: color = 2'b10;
      13'h10f6: color = 2'b11;
      13'h10f7: color = 2'b11;
      13'h10f8: color = 2'b10;
      13'h10f9: color = 2'b10;
      13'h10fa: color = 2'b11;
      13'h10fb: color = 2'b11;
      13'h10fc: color = 2'b11;
      13'h10fd: color = 2'b11;
      13'h10fe: color = 2'b11;
      13'h10ff: color = 2'b11;
      13'h1100: color = 2'b11;
      13'h1101: color = 2'b11;
      13'h1102: color = 2'b10;
      13'h1103: color = 2'b10;
      13'h1104: color = 2'b11;
      13'h1105: color = 2'b11;
      13'h1106: color = 2'b11;
      13'h1107: color = 2'b11;
      13'h1108: color = 2'b11;
      13'h1109: color = 2'b11;
      13'h110a: color = 2'b10;
      13'h110b: color = 2'b10;
      13'h110c: color = 2'b11;
      13'h110d: color = 2'b11;
      13'h110e: color = 2'b11;
      13'h110f: color = 2'b11;
      13'h1110: color = 2'b11;
      13'h1111: color = 2'b11;
      13'h1112: color = 2'b10;
      13'h1113: color = 2'b10;
      13'h1114: color = 2'b11;
      13'h1115: color = 2'b11;
      13'h1116: color = 2'b11;
      13'h1117: color = 2'b11;
      13'h1118: color = 2'b11;
      13'h1119: color = 2'b11;
      13'h111a: color = 2'b10;
      13'h111b: color = 2'b10;
      13'h111c: color = 2'b11;
      13'h111d: color = 2'b11;
      13'h111e: color = 2'b11;
      13'h111f: color = 2'b11;
      13'h1120: color = 2'b00;
      13'h1121: color = 2'b00;
      13'h1122: color = 2'b11;
      13'h1123: color = 2'b11;
      13'h1124: color = 2'b10;
      13'h1125: color = 2'b10;
      13'h1126: color = 2'b10;
      13'h1127: color = 2'b10;
      13'h1128: color = 2'b10;
      13'h1129: color = 2'b10;
      13'h112a: color = 2'b10;
      13'h112b: color = 2'b10;
      13'h112c: color = 2'b10;
      13'h112d: color = 2'b10;
      13'h112e: color = 2'b10;
      13'h112f: color = 2'b10;
      13'h1130: color = 2'b10;
      13'h1131: color = 2'b10;
      13'h1132: color = 2'b10;
      13'h1133: color = 2'b10;
      13'h1134: color = 2'b10;
      13'h1135: color = 2'b10;
      13'h1136: color = 2'b10;
      13'h1137: color = 2'b10;
      13'h1138: color = 2'b10;
      13'h1139: color = 2'b10;
      13'h113a: color = 2'b10;
      13'h113b: color = 2'b10;
      13'h113c: color = 2'b10;
      13'h113d: color = 2'b10;
      13'h113e: color = 2'b10;
      13'h113f: color = 2'b10;
      13'h1140: color = 2'b10;
      13'h1141: color = 2'b10;
      13'h1142: color = 2'b10;
      13'h1143: color = 2'b10;
      13'h1144: color = 2'b10;
      13'h1145: color = 2'b10;
      13'h1146: color = 2'b10;
      13'h1147: color = 2'b10;
      13'h1148: color = 2'b10;
      13'h1149: color = 2'b10;
      13'h114a: color = 2'b10;
      13'h114b: color = 2'b10;
      13'h114c: color = 2'b10;
      13'h114d: color = 2'b10;
      13'h114e: color = 2'b10;
      13'h114f: color = 2'b10;
      13'h1150: color = 2'b10;
      13'h1151: color = 2'b10;
      13'h1152: color = 2'b10;
      13'h1153: color = 2'b10;
      13'h1154: color = 2'b10;
      13'h1155: color = 2'b10;
      13'h1156: color = 2'b10;
      13'h1157: color = 2'b10;
      13'h1158: color = 2'b10;
      13'h1159: color = 2'b10;
      13'h115a: color = 2'b10;
      13'h115b: color = 2'b10;
      13'h115c: color = 2'b01;
      13'h115d: color = 2'b01;
      13'h115e: color = 2'b00;
      13'h115f: color = 2'b00;
      13'h1160: color = 2'b11;
      13'h1161: color = 2'b11;
      13'h1162: color = 2'b10;
      13'h1163: color = 2'b10;
      13'h1164: color = 2'b11;
      13'h1165: color = 2'b11;
      13'h1166: color = 2'b11;
      13'h1167: color = 2'b11;
      13'h1168: color = 2'b11;
      13'h1169: color = 2'b11;
      13'h116a: color = 2'b10;
      13'h116b: color = 2'b10;
      13'h116c: color = 2'b11;
      13'h116d: color = 2'b11;
      13'h116e: color = 2'b11;
      13'h116f: color = 2'b11;
      13'h1170: color = 2'b11;
      13'h1171: color = 2'b11;
      13'h1172: color = 2'b10;
      13'h1173: color = 2'b10;
      13'h1174: color = 2'b11;
      13'h1175: color = 2'b11;
      13'h1176: color = 2'b11;
      13'h1177: color = 2'b11;
      13'h1178: color = 2'b11;
      13'h1179: color = 2'b11;
      13'h117a: color = 2'b10;
      13'h117b: color = 2'b10;
      13'h117c: color = 2'b11;
      13'h117d: color = 2'b11;
      13'h117e: color = 2'b11;
      13'h117f: color = 2'b11;
      13'h1180: color = 2'b11;
      13'h1181: color = 2'b11;
      13'h1182: color = 2'b10;
      13'h1183: color = 2'b10;
      13'h1184: color = 2'b11;
      13'h1185: color = 2'b11;
      13'h1186: color = 2'b11;
      13'h1187: color = 2'b11;
      13'h1188: color = 2'b11;
      13'h1189: color = 2'b11;
      13'h118a: color = 2'b10;
      13'h118b: color = 2'b10;
      13'h118c: color = 2'b11;
      13'h118d: color = 2'b11;
      13'h118e: color = 2'b11;
      13'h118f: color = 2'b11;
      13'h1190: color = 2'b11;
      13'h1191: color = 2'b11;
      13'h1192: color = 2'b10;
      13'h1193: color = 2'b10;
      13'h1194: color = 2'b11;
      13'h1195: color = 2'b11;
      13'h1196: color = 2'b11;
      13'h1197: color = 2'b11;
      13'h1198: color = 2'b11;
      13'h1199: color = 2'b11;
      13'h119a: color = 2'b10;
      13'h119b: color = 2'b10;
      13'h119c: color = 2'b11;
      13'h119d: color = 2'b11;
      13'h119e: color = 2'b11;
      13'h119f: color = 2'b11;
      13'h11a0: color = 2'b00;
      13'h11a1: color = 2'b00;
      13'h11a2: color = 2'b11;
      13'h11a3: color = 2'b11;
      13'h11a4: color = 2'b10;
      13'h11a5: color = 2'b10;
      13'h11a6: color = 2'b10;
      13'h11a7: color = 2'b10;
      13'h11a8: color = 2'b10;
      13'h11a9: color = 2'b10;
      13'h11aa: color = 2'b10;
      13'h11ab: color = 2'b10;
      13'h11ac: color = 2'b10;
      13'h11ad: color = 2'b10;
      13'h11ae: color = 2'b10;
      13'h11af: color = 2'b10;
      13'h11b0: color = 2'b10;
      13'h11b1: color = 2'b10;
      13'h11b2: color = 2'b10;
      13'h11b3: color = 2'b10;
      13'h11b4: color = 2'b10;
      13'h11b5: color = 2'b10;
      13'h11b6: color = 2'b10;
      13'h11b7: color = 2'b10;
      13'h11b8: color = 2'b10;
      13'h11b9: color = 2'b10;
      13'h11ba: color = 2'b10;
      13'h11bb: color = 2'b10;
      13'h11bc: color = 2'b10;
      13'h11bd: color = 2'b10;
      13'h11be: color = 2'b10;
      13'h11bf: color = 2'b10;
      13'h11c0: color = 2'b10;
      13'h11c1: color = 2'b10;
      13'h11c2: color = 2'b10;
      13'h11c3: color = 2'b10;
      13'h11c4: color = 2'b10;
      13'h11c5: color = 2'b10;
      13'h11c6: color = 2'b10;
      13'h11c7: color = 2'b10;
      13'h11c8: color = 2'b10;
      13'h11c9: color = 2'b10;
      13'h11ca: color = 2'b10;
      13'h11cb: color = 2'b10;
      13'h11cc: color = 2'b10;
      13'h11cd: color = 2'b10;
      13'h11ce: color = 2'b10;
      13'h11cf: color = 2'b10;
      13'h11d0: color = 2'b10;
      13'h11d1: color = 2'b10;
      13'h11d2: color = 2'b10;
      13'h11d3: color = 2'b10;
      13'h11d4: color = 2'b10;
      13'h11d5: color = 2'b10;
      13'h11d6: color = 2'b10;
      13'h11d7: color = 2'b10;
      13'h11d8: color = 2'b10;
      13'h11d9: color = 2'b10;
      13'h11da: color = 2'b10;
      13'h11db: color = 2'b10;
      13'h11dc: color = 2'b01;
      13'h11dd: color = 2'b01;
      13'h11de: color = 2'b00;
      13'h11df: color = 2'b00;
      13'h11e0: color = 2'b11;
      13'h11e1: color = 2'b11;
      13'h11e2: color = 2'b10;
      13'h11e3: color = 2'b10;
      13'h11e4: color = 2'b11;
      13'h11e5: color = 2'b11;
      13'h11e6: color = 2'b11;
      13'h11e7: color = 2'b11;
      13'h11e8: color = 2'b11;
      13'h11e9: color = 2'b11;
      13'h11ea: color = 2'b10;
      13'h11eb: color = 2'b10;
      13'h11ec: color = 2'b11;
      13'h11ed: color = 2'b11;
      13'h11ee: color = 2'b11;
      13'h11ef: color = 2'b11;
      13'h11f0: color = 2'b11;
      13'h11f1: color = 2'b11;
      13'h11f2: color = 2'b10;
      13'h11f3: color = 2'b10;
      13'h11f4: color = 2'b11;
      13'h11f5: color = 2'b11;
      13'h11f6: color = 2'b11;
      13'h11f7: color = 2'b11;
      13'h11f8: color = 2'b11;
      13'h11f9: color = 2'b11;
      13'h11fa: color = 2'b10;
      13'h11fb: color = 2'b10;
      13'h11fc: color = 2'b11;
      13'h11fd: color = 2'b11;
      13'h11fe: color = 2'b11;
      13'h11ff: color = 2'b11;
      13'h1200: color = 2'b10;
      13'h1201: color = 2'b10;
      13'h1202: color = 2'b11;
      13'h1203: color = 2'b11;
      13'h1204: color = 2'b11;
      13'h1205: color = 2'b11;
      13'h1206: color = 2'b11;
      13'h1207: color = 2'b11;
      13'h1208: color = 2'b11;
      13'h1209: color = 2'b11;
      13'h120a: color = 2'b11;
      13'h120b: color = 2'b11;
      13'h120c: color = 2'b10;
      13'h120d: color = 2'b10;
      13'h120e: color = 2'b11;
      13'h120f: color = 2'b11;
      13'h1210: color = 2'b10;
      13'h1211: color = 2'b10;
      13'h1212: color = 2'b11;
      13'h1213: color = 2'b11;
      13'h1214: color = 2'b11;
      13'h1215: color = 2'b11;
      13'h1216: color = 2'b11;
      13'h1217: color = 2'b11;
      13'h1218: color = 2'b11;
      13'h1219: color = 2'b11;
      13'h121a: color = 2'b11;
      13'h121b: color = 2'b11;
      13'h121c: color = 2'b10;
      13'h121d: color = 2'b10;
      13'h121e: color = 2'b11;
      13'h121f: color = 2'b11;
      13'h1220: color = 2'b00;
      13'h1221: color = 2'b00;
      13'h1222: color = 2'b11;
      13'h1223: color = 2'b11;
      13'h1224: color = 2'b10;
      13'h1225: color = 2'b10;
      13'h1226: color = 2'b10;
      13'h1227: color = 2'b10;
      13'h1228: color = 2'b10;
      13'h1229: color = 2'b10;
      13'h122a: color = 2'b10;
      13'h122b: color = 2'b10;
      13'h122c: color = 2'b10;
      13'h122d: color = 2'b10;
      13'h122e: color = 2'b10;
      13'h122f: color = 2'b10;
      13'h1230: color = 2'b10;
      13'h1231: color = 2'b10;
      13'h1232: color = 2'b10;
      13'h1233: color = 2'b10;
      13'h1234: color = 2'b10;
      13'h1235: color = 2'b10;
      13'h1236: color = 2'b10;
      13'h1237: color = 2'b10;
      13'h1238: color = 2'b10;
      13'h1239: color = 2'b10;
      13'h123a: color = 2'b10;
      13'h123b: color = 2'b10;
      13'h123c: color = 2'b10;
      13'h123d: color = 2'b10;
      13'h123e: color = 2'b10;
      13'h123f: color = 2'b10;
      13'h1240: color = 2'b10;
      13'h1241: color = 2'b10;
      13'h1242: color = 2'b10;
      13'h1243: color = 2'b10;
      13'h1244: color = 2'b10;
      13'h1245: color = 2'b10;
      13'h1246: color = 2'b10;
      13'h1247: color = 2'b10;
      13'h1248: color = 2'b10;
      13'h1249: color = 2'b10;
      13'h124a: color = 2'b10;
      13'h124b: color = 2'b10;
      13'h124c: color = 2'b10;
      13'h124d: color = 2'b10;
      13'h124e: color = 2'b10;
      13'h124f: color = 2'b10;
      13'h1250: color = 2'b10;
      13'h1251: color = 2'b10;
      13'h1252: color = 2'b10;
      13'h1253: color = 2'b10;
      13'h1254: color = 2'b10;
      13'h1255: color = 2'b10;
      13'h1256: color = 2'b10;
      13'h1257: color = 2'b10;
      13'h1258: color = 2'b10;
      13'h1259: color = 2'b10;
      13'h125a: color = 2'b10;
      13'h125b: color = 2'b10;
      13'h125c: color = 2'b01;
      13'h125d: color = 2'b01;
      13'h125e: color = 2'b00;
      13'h125f: color = 2'b00;
      13'h1260: color = 2'b10;
      13'h1261: color = 2'b10;
      13'h1262: color = 2'b11;
      13'h1263: color = 2'b11;
      13'h1264: color = 2'b11;
      13'h1265: color = 2'b11;
      13'h1266: color = 2'b11;
      13'h1267: color = 2'b11;
      13'h1268: color = 2'b11;
      13'h1269: color = 2'b11;
      13'h126a: color = 2'b11;
      13'h126b: color = 2'b11;
      13'h126c: color = 2'b10;
      13'h126d: color = 2'b10;
      13'h126e: color = 2'b11;
      13'h126f: color = 2'b11;
      13'h1270: color = 2'b10;
      13'h1271: color = 2'b10;
      13'h1272: color = 2'b11;
      13'h1273: color = 2'b11;
      13'h1274: color = 2'b11;
      13'h1275: color = 2'b11;
      13'h1276: color = 2'b11;
      13'h1277: color = 2'b11;
      13'h1278: color = 2'b11;
      13'h1279: color = 2'b11;
      13'h127a: color = 2'b11;
      13'h127b: color = 2'b11;
      13'h127c: color = 2'b10;
      13'h127d: color = 2'b10;
      13'h127e: color = 2'b11;
      13'h127f: color = 2'b11;
      13'h1280: color = 2'b10;
      13'h1281: color = 2'b10;
      13'h1282: color = 2'b11;
      13'h1283: color = 2'b11;
      13'h1284: color = 2'b11;
      13'h1285: color = 2'b11;
      13'h1286: color = 2'b11;
      13'h1287: color = 2'b11;
      13'h1288: color = 2'b11;
      13'h1289: color = 2'b11;
      13'h128a: color = 2'b11;
      13'h128b: color = 2'b11;
      13'h128c: color = 2'b10;
      13'h128d: color = 2'b10;
      13'h128e: color = 2'b11;
      13'h128f: color = 2'b11;
      13'h1290: color = 2'b10;
      13'h1291: color = 2'b10;
      13'h1292: color = 2'b11;
      13'h1293: color = 2'b11;
      13'h1294: color = 2'b11;
      13'h1295: color = 2'b11;
      13'h1296: color = 2'b11;
      13'h1297: color = 2'b11;
      13'h1298: color = 2'b11;
      13'h1299: color = 2'b11;
      13'h129a: color = 2'b11;
      13'h129b: color = 2'b11;
      13'h129c: color = 2'b10;
      13'h129d: color = 2'b10;
      13'h129e: color = 2'b11;
      13'h129f: color = 2'b11;
      13'h12a0: color = 2'b00;
      13'h12a1: color = 2'b00;
      13'h12a2: color = 2'b11;
      13'h12a3: color = 2'b11;
      13'h12a4: color = 2'b10;
      13'h12a5: color = 2'b10;
      13'h12a6: color = 2'b10;
      13'h12a7: color = 2'b10;
      13'h12a8: color = 2'b10;
      13'h12a9: color = 2'b10;
      13'h12aa: color = 2'b10;
      13'h12ab: color = 2'b10;
      13'h12ac: color = 2'b10;
      13'h12ad: color = 2'b10;
      13'h12ae: color = 2'b10;
      13'h12af: color = 2'b10;
      13'h12b0: color = 2'b10;
      13'h12b1: color = 2'b10;
      13'h12b2: color = 2'b10;
      13'h12b3: color = 2'b10;
      13'h12b4: color = 2'b10;
      13'h12b5: color = 2'b10;
      13'h12b6: color = 2'b10;
      13'h12b7: color = 2'b10;
      13'h12b8: color = 2'b10;
      13'h12b9: color = 2'b10;
      13'h12ba: color = 2'b10;
      13'h12bb: color = 2'b10;
      13'h12bc: color = 2'b10;
      13'h12bd: color = 2'b10;
      13'h12be: color = 2'b10;
      13'h12bf: color = 2'b10;
      13'h12c0: color = 2'b10;
      13'h12c1: color = 2'b10;
      13'h12c2: color = 2'b10;
      13'h12c3: color = 2'b10;
      13'h12c4: color = 2'b10;
      13'h12c5: color = 2'b10;
      13'h12c6: color = 2'b10;
      13'h12c7: color = 2'b10;
      13'h12c8: color = 2'b10;
      13'h12c9: color = 2'b10;
      13'h12ca: color = 2'b10;
      13'h12cb: color = 2'b10;
      13'h12cc: color = 2'b10;
      13'h12cd: color = 2'b10;
      13'h12ce: color = 2'b10;
      13'h12cf: color = 2'b10;
      13'h12d0: color = 2'b10;
      13'h12d1: color = 2'b10;
      13'h12d2: color = 2'b10;
      13'h12d3: color = 2'b10;
      13'h12d4: color = 2'b10;
      13'h12d5: color = 2'b10;
      13'h12d6: color = 2'b10;
      13'h12d7: color = 2'b10;
      13'h12d8: color = 2'b10;
      13'h12d9: color = 2'b10;
      13'h12da: color = 2'b10;
      13'h12db: color = 2'b10;
      13'h12dc: color = 2'b01;
      13'h12dd: color = 2'b01;
      13'h12de: color = 2'b00;
      13'h12df: color = 2'b00;
      13'h12e0: color = 2'b10;
      13'h12e1: color = 2'b10;
      13'h12e2: color = 2'b11;
      13'h12e3: color = 2'b11;
      13'h12e4: color = 2'b11;
      13'h12e5: color = 2'b11;
      13'h12e6: color = 2'b11;
      13'h12e7: color = 2'b11;
      13'h12e8: color = 2'b11;
      13'h12e9: color = 2'b11;
      13'h12ea: color = 2'b11;
      13'h12eb: color = 2'b11;
      13'h12ec: color = 2'b10;
      13'h12ed: color = 2'b10;
      13'h12ee: color = 2'b11;
      13'h12ef: color = 2'b11;
      13'h12f0: color = 2'b10;
      13'h12f1: color = 2'b10;
      13'h12f2: color = 2'b11;
      13'h12f3: color = 2'b11;
      13'h12f4: color = 2'b11;
      13'h12f5: color = 2'b11;
      13'h12f6: color = 2'b11;
      13'h12f7: color = 2'b11;
      13'h12f8: color = 2'b11;
      13'h12f9: color = 2'b11;
      13'h12fa: color = 2'b11;
      13'h12fb: color = 2'b11;
      13'h12fc: color = 2'b10;
      13'h12fd: color = 2'b10;
      13'h12fe: color = 2'b11;
      13'h12ff: color = 2'b11;
      13'h1300: color = 2'b11;
      13'h1301: color = 2'b11;
      13'h1302: color = 2'b11;
      13'h1303: color = 2'b11;
      13'h1304: color = 2'b11;
      13'h1305: color = 2'b11;
      13'h1306: color = 2'b11;
      13'h1307: color = 2'b11;
      13'h1308: color = 2'b11;
      13'h1309: color = 2'b11;
      13'h130a: color = 2'b11;
      13'h130b: color = 2'b11;
      13'h130c: color = 2'b11;
      13'h130d: color = 2'b11;
      13'h130e: color = 2'b10;
      13'h130f: color = 2'b10;
      13'h1310: color = 2'b11;
      13'h1311: color = 2'b11;
      13'h1312: color = 2'b11;
      13'h1313: color = 2'b11;
      13'h1314: color = 2'b11;
      13'h1315: color = 2'b11;
      13'h1316: color = 2'b11;
      13'h1317: color = 2'b11;
      13'h1318: color = 2'b11;
      13'h1319: color = 2'b11;
      13'h131a: color = 2'b11;
      13'h131b: color = 2'b11;
      13'h131c: color = 2'b11;
      13'h131d: color = 2'b11;
      13'h131e: color = 2'b10;
      13'h131f: color = 2'b10;
      13'h1320: color = 2'b00;
      13'h1321: color = 2'b00;
      13'h1322: color = 2'b11;
      13'h1323: color = 2'b11;
      13'h1324: color = 2'b10;
      13'h1325: color = 2'b10;
      13'h1326: color = 2'b10;
      13'h1327: color = 2'b10;
      13'h1328: color = 2'b10;
      13'h1329: color = 2'b10;
      13'h132a: color = 2'b10;
      13'h132b: color = 2'b10;
      13'h132c: color = 2'b10;
      13'h132d: color = 2'b10;
      13'h132e: color = 2'b10;
      13'h132f: color = 2'b10;
      13'h1330: color = 2'b10;
      13'h1331: color = 2'b10;
      13'h1332: color = 2'b10;
      13'h1333: color = 2'b10;
      13'h1334: color = 2'b10;
      13'h1335: color = 2'b10;
      13'h1336: color = 2'b10;
      13'h1337: color = 2'b10;
      13'h1338: color = 2'b10;
      13'h1339: color = 2'b10;
      13'h133a: color = 2'b10;
      13'h133b: color = 2'b10;
      13'h133c: color = 2'b10;
      13'h133d: color = 2'b10;
      13'h133e: color = 2'b10;
      13'h133f: color = 2'b10;
      13'h1340: color = 2'b10;
      13'h1341: color = 2'b10;
      13'h1342: color = 2'b10;
      13'h1343: color = 2'b10;
      13'h1344: color = 2'b10;
      13'h1345: color = 2'b10;
      13'h1346: color = 2'b10;
      13'h1347: color = 2'b10;
      13'h1348: color = 2'b10;
      13'h1349: color = 2'b10;
      13'h134a: color = 2'b10;
      13'h134b: color = 2'b10;
      13'h134c: color = 2'b10;
      13'h134d: color = 2'b10;
      13'h134e: color = 2'b10;
      13'h134f: color = 2'b10;
      13'h1350: color = 2'b10;
      13'h1351: color = 2'b10;
      13'h1352: color = 2'b10;
      13'h1353: color = 2'b10;
      13'h1354: color = 2'b10;
      13'h1355: color = 2'b10;
      13'h1356: color = 2'b10;
      13'h1357: color = 2'b10;
      13'h1358: color = 2'b10;
      13'h1359: color = 2'b10;
      13'h135a: color = 2'b10;
      13'h135b: color = 2'b10;
      13'h135c: color = 2'b01;
      13'h135d: color = 2'b01;
      13'h135e: color = 2'b00;
      13'h135f: color = 2'b00;
      13'h1360: color = 2'b11;
      13'h1361: color = 2'b11;
      13'h1362: color = 2'b11;
      13'h1363: color = 2'b11;
      13'h1364: color = 2'b11;
      13'h1365: color = 2'b11;
      13'h1366: color = 2'b11;
      13'h1367: color = 2'b11;
      13'h1368: color = 2'b11;
      13'h1369: color = 2'b11;
      13'h136a: color = 2'b11;
      13'h136b: color = 2'b11;
      13'h136c: color = 2'b11;
      13'h136d: color = 2'b11;
      13'h136e: color = 2'b10;
      13'h136f: color = 2'b10;
      13'h1370: color = 2'b11;
      13'h1371: color = 2'b11;
      13'h1372: color = 2'b11;
      13'h1373: color = 2'b11;
      13'h1374: color = 2'b11;
      13'h1375: color = 2'b11;
      13'h1376: color = 2'b11;
      13'h1377: color = 2'b11;
      13'h1378: color = 2'b11;
      13'h1379: color = 2'b11;
      13'h137a: color = 2'b11;
      13'h137b: color = 2'b11;
      13'h137c: color = 2'b11;
      13'h137d: color = 2'b11;
      13'h137e: color = 2'b10;
      13'h137f: color = 2'b10;
      13'h1380: color = 2'b11;
      13'h1381: color = 2'b11;
      13'h1382: color = 2'b11;
      13'h1383: color = 2'b11;
      13'h1384: color = 2'b11;
      13'h1385: color = 2'b11;
      13'h1386: color = 2'b11;
      13'h1387: color = 2'b11;
      13'h1388: color = 2'b11;
      13'h1389: color = 2'b11;
      13'h138a: color = 2'b11;
      13'h138b: color = 2'b11;
      13'h138c: color = 2'b11;
      13'h138d: color = 2'b11;
      13'h138e: color = 2'b10;
      13'h138f: color = 2'b10;
      13'h1390: color = 2'b11;
      13'h1391: color = 2'b11;
      13'h1392: color = 2'b11;
      13'h1393: color = 2'b11;
      13'h1394: color = 2'b11;
      13'h1395: color = 2'b11;
      13'h1396: color = 2'b11;
      13'h1397: color = 2'b11;
      13'h1398: color = 2'b11;
      13'h1399: color = 2'b11;
      13'h139a: color = 2'b11;
      13'h139b: color = 2'b11;
      13'h139c: color = 2'b11;
      13'h139d: color = 2'b11;
      13'h139e: color = 2'b10;
      13'h139f: color = 2'b10;
      13'h13a0: color = 2'b00;
      13'h13a1: color = 2'b00;
      13'h13a2: color = 2'b11;
      13'h13a3: color = 2'b11;
      13'h13a4: color = 2'b10;
      13'h13a5: color = 2'b10;
      13'h13a6: color = 2'b10;
      13'h13a7: color = 2'b10;
      13'h13a8: color = 2'b10;
      13'h13a9: color = 2'b10;
      13'h13aa: color = 2'b10;
      13'h13ab: color = 2'b10;
      13'h13ac: color = 2'b10;
      13'h13ad: color = 2'b10;
      13'h13ae: color = 2'b10;
      13'h13af: color = 2'b10;
      13'h13b0: color = 2'b10;
      13'h13b1: color = 2'b10;
      13'h13b2: color = 2'b10;
      13'h13b3: color = 2'b10;
      13'h13b4: color = 2'b10;
      13'h13b5: color = 2'b10;
      13'h13b6: color = 2'b10;
      13'h13b7: color = 2'b10;
      13'h13b8: color = 2'b10;
      13'h13b9: color = 2'b10;
      13'h13ba: color = 2'b10;
      13'h13bb: color = 2'b10;
      13'h13bc: color = 2'b10;
      13'h13bd: color = 2'b10;
      13'h13be: color = 2'b10;
      13'h13bf: color = 2'b10;
      13'h13c0: color = 2'b10;
      13'h13c1: color = 2'b10;
      13'h13c2: color = 2'b10;
      13'h13c3: color = 2'b10;
      13'h13c4: color = 2'b10;
      13'h13c5: color = 2'b10;
      13'h13c6: color = 2'b10;
      13'h13c7: color = 2'b10;
      13'h13c8: color = 2'b10;
      13'h13c9: color = 2'b10;
      13'h13ca: color = 2'b10;
      13'h13cb: color = 2'b10;
      13'h13cc: color = 2'b10;
      13'h13cd: color = 2'b10;
      13'h13ce: color = 2'b10;
      13'h13cf: color = 2'b10;
      13'h13d0: color = 2'b10;
      13'h13d1: color = 2'b10;
      13'h13d2: color = 2'b10;
      13'h13d3: color = 2'b10;
      13'h13d4: color = 2'b10;
      13'h13d5: color = 2'b10;
      13'h13d6: color = 2'b10;
      13'h13d7: color = 2'b10;
      13'h13d8: color = 2'b10;
      13'h13d9: color = 2'b10;
      13'h13da: color = 2'b10;
      13'h13db: color = 2'b10;
      13'h13dc: color = 2'b01;
      13'h13dd: color = 2'b01;
      13'h13de: color = 2'b00;
      13'h13df: color = 2'b00;
      13'h13e0: color = 2'b11;
      13'h13e1: color = 2'b11;
      13'h13e2: color = 2'b11;
      13'h13e3: color = 2'b11;
      13'h13e4: color = 2'b11;
      13'h13e5: color = 2'b11;
      13'h13e6: color = 2'b11;
      13'h13e7: color = 2'b11;
      13'h13e8: color = 2'b11;
      13'h13e9: color = 2'b11;
      13'h13ea: color = 2'b11;
      13'h13eb: color = 2'b11;
      13'h13ec: color = 2'b11;
      13'h13ed: color = 2'b11;
      13'h13ee: color = 2'b10;
      13'h13ef: color = 2'b10;
      13'h13f0: color = 2'b11;
      13'h13f1: color = 2'b11;
      13'h13f2: color = 2'b11;
      13'h13f3: color = 2'b11;
      13'h13f4: color = 2'b11;
      13'h13f5: color = 2'b11;
      13'h13f6: color = 2'b11;
      13'h13f7: color = 2'b11;
      13'h13f8: color = 2'b11;
      13'h13f9: color = 2'b11;
      13'h13fa: color = 2'b11;
      13'h13fb: color = 2'b11;
      13'h13fc: color = 2'b11;
      13'h13fd: color = 2'b11;
      13'h13fe: color = 2'b10;
      13'h13ff: color = 2'b10;
      13'h1400: color = 2'b10;
      13'h1401: color = 2'b10;
      13'h1402: color = 2'b11;
      13'h1403: color = 2'b11;
      13'h1404: color = 2'b11;
      13'h1405: color = 2'b11;
      13'h1406: color = 2'b11;
      13'h1407: color = 2'b11;
      13'h1408: color = 2'b11;
      13'h1409: color = 2'b11;
      13'h140a: color = 2'b11;
      13'h140b: color = 2'b11;
      13'h140c: color = 2'b11;
      13'h140d: color = 2'b11;
      13'h140e: color = 2'b11;
      13'h140f: color = 2'b11;
      13'h1410: color = 2'b10;
      13'h1411: color = 2'b10;
      13'h1412: color = 2'b11;
      13'h1413: color = 2'b11;
      13'h1414: color = 2'b11;
      13'h1415: color = 2'b11;
      13'h1416: color = 2'b11;
      13'h1417: color = 2'b11;
      13'h1418: color = 2'b11;
      13'h1419: color = 2'b11;
      13'h141a: color = 2'b11;
      13'h141b: color = 2'b11;
      13'h141c: color = 2'b11;
      13'h141d: color = 2'b11;
      13'h141e: color = 2'b11;
      13'h141f: color = 2'b11;
      13'h1420: color = 2'b00;
      13'h1421: color = 2'b00;
      13'h1422: color = 2'b11;
      13'h1423: color = 2'b11;
      13'h1424: color = 2'b10;
      13'h1425: color = 2'b10;
      13'h1426: color = 2'b10;
      13'h1427: color = 2'b10;
      13'h1428: color = 2'b10;
      13'h1429: color = 2'b10;
      13'h142a: color = 2'b10;
      13'h142b: color = 2'b10;
      13'h142c: color = 2'b10;
      13'h142d: color = 2'b10;
      13'h142e: color = 2'b10;
      13'h142f: color = 2'b10;
      13'h1430: color = 2'b10;
      13'h1431: color = 2'b10;
      13'h1432: color = 2'b10;
      13'h1433: color = 2'b10;
      13'h1434: color = 2'b10;
      13'h1435: color = 2'b10;
      13'h1436: color = 2'b10;
      13'h1437: color = 2'b10;
      13'h1438: color = 2'b10;
      13'h1439: color = 2'b10;
      13'h143a: color = 2'b10;
      13'h143b: color = 2'b10;
      13'h143c: color = 2'b10;
      13'h143d: color = 2'b10;
      13'h143e: color = 2'b10;
      13'h143f: color = 2'b10;
      13'h1440: color = 2'b10;
      13'h1441: color = 2'b10;
      13'h1442: color = 2'b10;
      13'h1443: color = 2'b10;
      13'h1444: color = 2'b10;
      13'h1445: color = 2'b10;
      13'h1446: color = 2'b10;
      13'h1447: color = 2'b10;
      13'h1448: color = 2'b10;
      13'h1449: color = 2'b10;
      13'h144a: color = 2'b10;
      13'h144b: color = 2'b10;
      13'h144c: color = 2'b10;
      13'h144d: color = 2'b10;
      13'h144e: color = 2'b10;
      13'h144f: color = 2'b10;
      13'h1450: color = 2'b10;
      13'h1451: color = 2'b10;
      13'h1452: color = 2'b10;
      13'h1453: color = 2'b10;
      13'h1454: color = 2'b10;
      13'h1455: color = 2'b10;
      13'h1456: color = 2'b10;
      13'h1457: color = 2'b10;
      13'h1458: color = 2'b10;
      13'h1459: color = 2'b10;
      13'h145a: color = 2'b10;
      13'h145b: color = 2'b10;
      13'h145c: color = 2'b01;
      13'h145d: color = 2'b01;
      13'h145e: color = 2'b00;
      13'h145f: color = 2'b00;
      13'h1460: color = 2'b10;
      13'h1461: color = 2'b10;
      13'h1462: color = 2'b11;
      13'h1463: color = 2'b11;
      13'h1464: color = 2'b11;
      13'h1465: color = 2'b11;
      13'h1466: color = 2'b11;
      13'h1467: color = 2'b11;
      13'h1468: color = 2'b11;
      13'h1469: color = 2'b11;
      13'h146a: color = 2'b11;
      13'h146b: color = 2'b11;
      13'h146c: color = 2'b11;
      13'h146d: color = 2'b11;
      13'h146e: color = 2'b11;
      13'h146f: color = 2'b11;
      13'h1470: color = 2'b10;
      13'h1471: color = 2'b10;
      13'h1472: color = 2'b11;
      13'h1473: color = 2'b11;
      13'h1474: color = 2'b11;
      13'h1475: color = 2'b11;
      13'h1476: color = 2'b11;
      13'h1477: color = 2'b11;
      13'h1478: color = 2'b11;
      13'h1479: color = 2'b11;
      13'h147a: color = 2'b11;
      13'h147b: color = 2'b11;
      13'h147c: color = 2'b11;
      13'h147d: color = 2'b11;
      13'h147e: color = 2'b11;
      13'h147f: color = 2'b11;
      13'h1480: color = 2'b10;
      13'h1481: color = 2'b10;
      13'h1482: color = 2'b11;
      13'h1483: color = 2'b11;
      13'h1484: color = 2'b11;
      13'h1485: color = 2'b11;
      13'h1486: color = 2'b11;
      13'h1487: color = 2'b11;
      13'h1488: color = 2'b11;
      13'h1489: color = 2'b11;
      13'h148a: color = 2'b11;
      13'h148b: color = 2'b11;
      13'h148c: color = 2'b11;
      13'h148d: color = 2'b11;
      13'h148e: color = 2'b11;
      13'h148f: color = 2'b11;
      13'h1490: color = 2'b10;
      13'h1491: color = 2'b10;
      13'h1492: color = 2'b11;
      13'h1493: color = 2'b11;
      13'h1494: color = 2'b11;
      13'h1495: color = 2'b11;
      13'h1496: color = 2'b11;
      13'h1497: color = 2'b11;
      13'h1498: color = 2'b11;
      13'h1499: color = 2'b11;
      13'h149a: color = 2'b11;
      13'h149b: color = 2'b11;
      13'h149c: color = 2'b11;
      13'h149d: color = 2'b11;
      13'h149e: color = 2'b11;
      13'h149f: color = 2'b11;
      13'h14a0: color = 2'b00;
      13'h14a1: color = 2'b00;
      13'h14a2: color = 2'b11;
      13'h14a3: color = 2'b11;
      13'h14a4: color = 2'b10;
      13'h14a5: color = 2'b10;
      13'h14a6: color = 2'b10;
      13'h14a7: color = 2'b10;
      13'h14a8: color = 2'b10;
      13'h14a9: color = 2'b10;
      13'h14aa: color = 2'b10;
      13'h14ab: color = 2'b10;
      13'h14ac: color = 2'b10;
      13'h14ad: color = 2'b10;
      13'h14ae: color = 2'b10;
      13'h14af: color = 2'b10;
      13'h14b0: color = 2'b10;
      13'h14b1: color = 2'b10;
      13'h14b2: color = 2'b10;
      13'h14b3: color = 2'b10;
      13'h14b4: color = 2'b10;
      13'h14b5: color = 2'b10;
      13'h14b6: color = 2'b10;
      13'h14b7: color = 2'b10;
      13'h14b8: color = 2'b10;
      13'h14b9: color = 2'b10;
      13'h14ba: color = 2'b10;
      13'h14bb: color = 2'b10;
      13'h14bc: color = 2'b10;
      13'h14bd: color = 2'b10;
      13'h14be: color = 2'b10;
      13'h14bf: color = 2'b10;
      13'h14c0: color = 2'b10;
      13'h14c1: color = 2'b10;
      13'h14c2: color = 2'b10;
      13'h14c3: color = 2'b10;
      13'h14c4: color = 2'b10;
      13'h14c5: color = 2'b10;
      13'h14c6: color = 2'b10;
      13'h14c7: color = 2'b10;
      13'h14c8: color = 2'b10;
      13'h14c9: color = 2'b10;
      13'h14ca: color = 2'b10;
      13'h14cb: color = 2'b10;
      13'h14cc: color = 2'b10;
      13'h14cd: color = 2'b10;
      13'h14ce: color = 2'b10;
      13'h14cf: color = 2'b10;
      13'h14d0: color = 2'b10;
      13'h14d1: color = 2'b10;
      13'h14d2: color = 2'b10;
      13'h14d3: color = 2'b10;
      13'h14d4: color = 2'b10;
      13'h14d5: color = 2'b10;
      13'h14d6: color = 2'b10;
      13'h14d7: color = 2'b10;
      13'h14d8: color = 2'b10;
      13'h14d9: color = 2'b10;
      13'h14da: color = 2'b10;
      13'h14db: color = 2'b10;
      13'h14dc: color = 2'b01;
      13'h14dd: color = 2'b01;
      13'h14de: color = 2'b00;
      13'h14df: color = 2'b00;
      13'h14e0: color = 2'b10;
      13'h14e1: color = 2'b10;
      13'h14e2: color = 2'b11;
      13'h14e3: color = 2'b11;
      13'h14e4: color = 2'b11;
      13'h14e5: color = 2'b11;
      13'h14e6: color = 2'b11;
      13'h14e7: color = 2'b11;
      13'h14e8: color = 2'b11;
      13'h14e9: color = 2'b11;
      13'h14ea: color = 2'b11;
      13'h14eb: color = 2'b11;
      13'h14ec: color = 2'b11;
      13'h14ed: color = 2'b11;
      13'h14ee: color = 2'b11;
      13'h14ef: color = 2'b11;
      13'h14f0: color = 2'b10;
      13'h14f1: color = 2'b10;
      13'h14f2: color = 2'b11;
      13'h14f3: color = 2'b11;
      13'h14f4: color = 2'b11;
      13'h14f5: color = 2'b11;
      13'h14f6: color = 2'b11;
      13'h14f7: color = 2'b11;
      13'h14f8: color = 2'b11;
      13'h14f9: color = 2'b11;
      13'h14fa: color = 2'b11;
      13'h14fb: color = 2'b11;
      13'h14fc: color = 2'b11;
      13'h14fd: color = 2'b11;
      13'h14fe: color = 2'b11;
      13'h14ff: color = 2'b11;
      13'h1500: color = 2'b11;
      13'h1501: color = 2'b11;
      13'h1502: color = 2'b10;
      13'h1503: color = 2'b10;
      13'h1504: color = 2'b11;
      13'h1505: color = 2'b11;
      13'h1506: color = 2'b00;
      13'h1507: color = 2'b00;
      13'h1508: color = 2'b00;
      13'h1509: color = 2'b00;
      13'h150a: color = 2'b00;
      13'h150b: color = 2'b00;
      13'h150c: color = 2'b00;
      13'h150d: color = 2'b00;
      13'h150e: color = 2'b00;
      13'h150f: color = 2'b00;
      13'h1510: color = 2'b00;
      13'h1511: color = 2'b00;
      13'h1512: color = 2'b00;
      13'h1513: color = 2'b00;
      13'h1514: color = 2'b00;
      13'h1515: color = 2'b00;
      13'h1516: color = 2'b00;
      13'h1517: color = 2'b00;
      13'h1518: color = 2'b00;
      13'h1519: color = 2'b00;
      13'h151a: color = 2'b11;
      13'h151b: color = 2'b11;
      13'h151c: color = 2'b11;
      13'h151d: color = 2'b11;
      13'h151e: color = 2'b11;
      13'h151f: color = 2'b11;
      13'h1520: color = 2'b00;
      13'h1521: color = 2'b00;
      13'h1522: color = 2'b11;
      13'h1523: color = 2'b11;
      13'h1524: color = 2'b10;
      13'h1525: color = 2'b10;
      13'h1526: color = 2'b10;
      13'h1527: color = 2'b10;
      13'h1528: color = 2'b10;
      13'h1529: color = 2'b10;
      13'h152a: color = 2'b10;
      13'h152b: color = 2'b10;
      13'h152c: color = 2'b10;
      13'h152d: color = 2'b10;
      13'h152e: color = 2'b10;
      13'h152f: color = 2'b10;
      13'h1530: color = 2'b10;
      13'h1531: color = 2'b10;
      13'h1532: color = 2'b10;
      13'h1533: color = 2'b10;
      13'h1534: color = 2'b10;
      13'h1535: color = 2'b10;
      13'h1536: color = 2'b10;
      13'h1537: color = 2'b10;
      13'h1538: color = 2'b10;
      13'h1539: color = 2'b10;
      13'h153a: color = 2'b10;
      13'h153b: color = 2'b10;
      13'h153c: color = 2'b10;
      13'h153d: color = 2'b10;
      13'h153e: color = 2'b10;
      13'h153f: color = 2'b10;
      13'h1540: color = 2'b10;
      13'h1541: color = 2'b10;
      13'h1542: color = 2'b10;
      13'h1543: color = 2'b10;
      13'h1544: color = 2'b10;
      13'h1545: color = 2'b10;
      13'h1546: color = 2'b10;
      13'h1547: color = 2'b10;
      13'h1548: color = 2'b10;
      13'h1549: color = 2'b10;
      13'h154a: color = 2'b10;
      13'h154b: color = 2'b10;
      13'h154c: color = 2'b10;
      13'h154d: color = 2'b10;
      13'h154e: color = 2'b10;
      13'h154f: color = 2'b10;
      13'h1550: color = 2'b10;
      13'h1551: color = 2'b10;
      13'h1552: color = 2'b10;
      13'h1553: color = 2'b10;
      13'h1554: color = 2'b10;
      13'h1555: color = 2'b10;
      13'h1556: color = 2'b10;
      13'h1557: color = 2'b10;
      13'h1558: color = 2'b10;
      13'h1559: color = 2'b10;
      13'h155a: color = 2'b10;
      13'h155b: color = 2'b10;
      13'h155c: color = 2'b01;
      13'h155d: color = 2'b01;
      13'h155e: color = 2'b00;
      13'h155f: color = 2'b00;
      13'h1560: color = 2'b11;
      13'h1561: color = 2'b11;
      13'h1562: color = 2'b10;
      13'h1563: color = 2'b10;
      13'h1564: color = 2'b11;
      13'h1565: color = 2'b11;
      13'h1566: color = 2'b00;
      13'h1567: color = 2'b00;
      13'h1568: color = 2'b00;
      13'h1569: color = 2'b00;
      13'h156a: color = 2'b00;
      13'h156b: color = 2'b00;
      13'h156c: color = 2'b00;
      13'h156d: color = 2'b00;
      13'h156e: color = 2'b00;
      13'h156f: color = 2'b00;
      13'h1570: color = 2'b00;
      13'h1571: color = 2'b00;
      13'h1572: color = 2'b00;
      13'h1573: color = 2'b00;
      13'h1574: color = 2'b00;
      13'h1575: color = 2'b00;
      13'h1576: color = 2'b00;
      13'h1577: color = 2'b00;
      13'h1578: color = 2'b00;
      13'h1579: color = 2'b00;
      13'h157a: color = 2'b11;
      13'h157b: color = 2'b11;
      13'h157c: color = 2'b11;
      13'h157d: color = 2'b11;
      13'h157e: color = 2'b11;
      13'h157f: color = 2'b11;
      13'h1580: color = 2'b11;
      13'h1581: color = 2'b11;
      13'h1582: color = 2'b10;
      13'h1583: color = 2'b10;
      13'h1584: color = 2'b11;
      13'h1585: color = 2'b11;
      13'h1586: color = 2'b00;
      13'h1587: color = 2'b00;
      13'h1588: color = 2'b00;
      13'h1589: color = 2'b00;
      13'h158a: color = 2'b00;
      13'h158b: color = 2'b00;
      13'h158c: color = 2'b00;
      13'h158d: color = 2'b00;
      13'h158e: color = 2'b00;
      13'h158f: color = 2'b00;
      13'h1590: color = 2'b00;
      13'h1591: color = 2'b00;
      13'h1592: color = 2'b00;
      13'h1593: color = 2'b00;
      13'h1594: color = 2'b00;
      13'h1595: color = 2'b00;
      13'h1596: color = 2'b00;
      13'h1597: color = 2'b00;
      13'h1598: color = 2'b00;
      13'h1599: color = 2'b00;
      13'h159a: color = 2'b11;
      13'h159b: color = 2'b11;
      13'h159c: color = 2'b11;
      13'h159d: color = 2'b11;
      13'h159e: color = 2'b11;
      13'h159f: color = 2'b11;
      13'h15a0: color = 2'b00;
      13'h15a1: color = 2'b00;
      13'h15a2: color = 2'b11;
      13'h15a3: color = 2'b11;
      13'h15a4: color = 2'b10;
      13'h15a5: color = 2'b10;
      13'h15a6: color = 2'b10;
      13'h15a7: color = 2'b10;
      13'h15a8: color = 2'b10;
      13'h15a9: color = 2'b10;
      13'h15aa: color = 2'b10;
      13'h15ab: color = 2'b10;
      13'h15ac: color = 2'b10;
      13'h15ad: color = 2'b10;
      13'h15ae: color = 2'b10;
      13'h15af: color = 2'b10;
      13'h15b0: color = 2'b10;
      13'h15b1: color = 2'b10;
      13'h15b2: color = 2'b10;
      13'h15b3: color = 2'b10;
      13'h15b4: color = 2'b10;
      13'h15b5: color = 2'b10;
      13'h15b6: color = 2'b10;
      13'h15b7: color = 2'b10;
      13'h15b8: color = 2'b10;
      13'h15b9: color = 2'b10;
      13'h15ba: color = 2'b10;
      13'h15bb: color = 2'b10;
      13'h15bc: color = 2'b10;
      13'h15bd: color = 2'b10;
      13'h15be: color = 2'b10;
      13'h15bf: color = 2'b10;
      13'h15c0: color = 2'b10;
      13'h15c1: color = 2'b10;
      13'h15c2: color = 2'b10;
      13'h15c3: color = 2'b10;
      13'h15c4: color = 2'b10;
      13'h15c5: color = 2'b10;
      13'h15c6: color = 2'b10;
      13'h15c7: color = 2'b10;
      13'h15c8: color = 2'b10;
      13'h15c9: color = 2'b10;
      13'h15ca: color = 2'b10;
      13'h15cb: color = 2'b10;
      13'h15cc: color = 2'b10;
      13'h15cd: color = 2'b10;
      13'h15ce: color = 2'b10;
      13'h15cf: color = 2'b10;
      13'h15d0: color = 2'b10;
      13'h15d1: color = 2'b10;
      13'h15d2: color = 2'b10;
      13'h15d3: color = 2'b10;
      13'h15d4: color = 2'b10;
      13'h15d5: color = 2'b10;
      13'h15d6: color = 2'b10;
      13'h15d7: color = 2'b10;
      13'h15d8: color = 2'b10;
      13'h15d9: color = 2'b10;
      13'h15da: color = 2'b10;
      13'h15db: color = 2'b10;
      13'h15dc: color = 2'b01;
      13'h15dd: color = 2'b01;
      13'h15de: color = 2'b00;
      13'h15df: color = 2'b00;
      13'h15e0: color = 2'b11;
      13'h15e1: color = 2'b11;
      13'h15e2: color = 2'b10;
      13'h15e3: color = 2'b10;
      13'h15e4: color = 2'b11;
      13'h15e5: color = 2'b11;
      13'h15e6: color = 2'b00;
      13'h15e7: color = 2'b00;
      13'h15e8: color = 2'b00;
      13'h15e9: color = 2'b00;
      13'h15ea: color = 2'b00;
      13'h15eb: color = 2'b00;
      13'h15ec: color = 2'b00;
      13'h15ed: color = 2'b00;
      13'h15ee: color = 2'b00;
      13'h15ef: color = 2'b00;
      13'h15f0: color = 2'b00;
      13'h15f1: color = 2'b00;
      13'h15f2: color = 2'b00;
      13'h15f3: color = 2'b00;
      13'h15f4: color = 2'b00;
      13'h15f5: color = 2'b00;
      13'h15f6: color = 2'b00;
      13'h15f7: color = 2'b00;
      13'h15f8: color = 2'b00;
      13'h15f9: color = 2'b00;
      13'h15fa: color = 2'b11;
      13'h15fb: color = 2'b11;
      13'h15fc: color = 2'b11;
      13'h15fd: color = 2'b11;
      13'h15fe: color = 2'b11;
      13'h15ff: color = 2'b11;
      13'h1600: color = 2'b11;
      13'h1601: color = 2'b11;
      13'h1602: color = 2'b11;
      13'h1603: color = 2'b11;
      13'h1604: color = 2'b00;
      13'h1605: color = 2'b00;
      13'h1606: color = 2'b11;
      13'h1607: color = 2'b11;
      13'h1608: color = 2'b11;
      13'h1609: color = 2'b11;
      13'h160a: color = 2'b11;
      13'h160b: color = 2'b11;
      13'h160c: color = 2'b11;
      13'h160d: color = 2'b11;
      13'h160e: color = 2'b11;
      13'h160f: color = 2'b11;
      13'h1610: color = 2'b11;
      13'h1611: color = 2'b11;
      13'h1612: color = 2'b11;
      13'h1613: color = 2'b11;
      13'h1614: color = 2'b11;
      13'h1615: color = 2'b11;
      13'h1616: color = 2'b11;
      13'h1617: color = 2'b11;
      13'h1618: color = 2'b11;
      13'h1619: color = 2'b11;
      13'h161a: color = 2'b00;
      13'h161b: color = 2'b00;
      13'h161c: color = 2'b11;
      13'h161d: color = 2'b11;
      13'h161e: color = 2'b11;
      13'h161f: color = 2'b11;
      13'h1620: color = 2'b00;
      13'h1621: color = 2'b00;
      13'h1622: color = 2'b11;
      13'h1623: color = 2'b11;
      13'h1624: color = 2'b10;
      13'h1625: color = 2'b10;
      13'h1626: color = 2'b10;
      13'h1627: color = 2'b10;
      13'h1628: color = 2'b10;
      13'h1629: color = 2'b10;
      13'h162a: color = 2'b10;
      13'h162b: color = 2'b10;
      13'h162c: color = 2'b10;
      13'h162d: color = 2'b10;
      13'h162e: color = 2'b10;
      13'h162f: color = 2'b10;
      13'h1630: color = 2'b10;
      13'h1631: color = 2'b10;
      13'h1632: color = 2'b10;
      13'h1633: color = 2'b10;
      13'h1634: color = 2'b10;
      13'h1635: color = 2'b10;
      13'h1636: color = 2'b10;
      13'h1637: color = 2'b10;
      13'h1638: color = 2'b10;
      13'h1639: color = 2'b10;
      13'h163a: color = 2'b10;
      13'h163b: color = 2'b10;
      13'h163c: color = 2'b10;
      13'h163d: color = 2'b10;
      13'h163e: color = 2'b10;
      13'h163f: color = 2'b10;
      13'h1640: color = 2'b10;
      13'h1641: color = 2'b10;
      13'h1642: color = 2'b10;
      13'h1643: color = 2'b10;
      13'h1644: color = 2'b10;
      13'h1645: color = 2'b10;
      13'h1646: color = 2'b10;
      13'h1647: color = 2'b10;
      13'h1648: color = 2'b10;
      13'h1649: color = 2'b10;
      13'h164a: color = 2'b10;
      13'h164b: color = 2'b10;
      13'h164c: color = 2'b10;
      13'h164d: color = 2'b10;
      13'h164e: color = 2'b10;
      13'h164f: color = 2'b10;
      13'h1650: color = 2'b10;
      13'h1651: color = 2'b10;
      13'h1652: color = 2'b10;
      13'h1653: color = 2'b10;
      13'h1654: color = 2'b10;
      13'h1655: color = 2'b10;
      13'h1656: color = 2'b10;
      13'h1657: color = 2'b10;
      13'h1658: color = 2'b10;
      13'h1659: color = 2'b10;
      13'h165a: color = 2'b10;
      13'h165b: color = 2'b10;
      13'h165c: color = 2'b01;
      13'h165d: color = 2'b01;
      13'h165e: color = 2'b00;
      13'h165f: color = 2'b00;
      13'h1660: color = 2'b11;
      13'h1661: color = 2'b11;
      13'h1662: color = 2'b11;
      13'h1663: color = 2'b11;
      13'h1664: color = 2'b00;
      13'h1665: color = 2'b00;
      13'h1666: color = 2'b11;
      13'h1667: color = 2'b11;
      13'h1668: color = 2'b11;
      13'h1669: color = 2'b11;
      13'h166a: color = 2'b11;
      13'h166b: color = 2'b11;
      13'h166c: color = 2'b11;
      13'h166d: color = 2'b11;
      13'h166e: color = 2'b11;
      13'h166f: color = 2'b11;
      13'h1670: color = 2'b11;
      13'h1671: color = 2'b11;
      13'h1672: color = 2'b11;
      13'h1673: color = 2'b11;
      13'h1674: color = 2'b11;
      13'h1675: color = 2'b11;
      13'h1676: color = 2'b11;
      13'h1677: color = 2'b11;
      13'h1678: color = 2'b11;
      13'h1679: color = 2'b11;
      13'h167a: color = 2'b00;
      13'h167b: color = 2'b00;
      13'h167c: color = 2'b11;
      13'h167d: color = 2'b11;
      13'h167e: color = 2'b11;
      13'h167f: color = 2'b11;
      13'h1680: color = 2'b11;
      13'h1681: color = 2'b11;
      13'h1682: color = 2'b11;
      13'h1683: color = 2'b11;
      13'h1684: color = 2'b00;
      13'h1685: color = 2'b00;
      13'h1686: color = 2'b11;
      13'h1687: color = 2'b11;
      13'h1688: color = 2'b11;
      13'h1689: color = 2'b11;
      13'h168a: color = 2'b11;
      13'h168b: color = 2'b11;
      13'h168c: color = 2'b11;
      13'h168d: color = 2'b11;
      13'h168e: color = 2'b11;
      13'h168f: color = 2'b11;
      13'h1690: color = 2'b11;
      13'h1691: color = 2'b11;
      13'h1692: color = 2'b11;
      13'h1693: color = 2'b11;
      13'h1694: color = 2'b11;
      13'h1695: color = 2'b11;
      13'h1696: color = 2'b11;
      13'h1697: color = 2'b11;
      13'h1698: color = 2'b11;
      13'h1699: color = 2'b11;
      13'h169a: color = 2'b00;
      13'h169b: color = 2'b00;
      13'h169c: color = 2'b11;
      13'h169d: color = 2'b11;
      13'h169e: color = 2'b11;
      13'h169f: color = 2'b11;
      13'h16a0: color = 2'b00;
      13'h16a1: color = 2'b00;
      13'h16a2: color = 2'b11;
      13'h16a3: color = 2'b11;
      13'h16a4: color = 2'b10;
      13'h16a5: color = 2'b10;
      13'h16a6: color = 2'b10;
      13'h16a7: color = 2'b10;
      13'h16a8: color = 2'b10;
      13'h16a9: color = 2'b10;
      13'h16aa: color = 2'b10;
      13'h16ab: color = 2'b10;
      13'h16ac: color = 2'b10;
      13'h16ad: color = 2'b10;
      13'h16ae: color = 2'b10;
      13'h16af: color = 2'b10;
      13'h16b0: color = 2'b10;
      13'h16b1: color = 2'b10;
      13'h16b2: color = 2'b10;
      13'h16b3: color = 2'b10;
      13'h16b4: color = 2'b10;
      13'h16b5: color = 2'b10;
      13'h16b6: color = 2'b10;
      13'h16b7: color = 2'b10;
      13'h16b8: color = 2'b10;
      13'h16b9: color = 2'b10;
      13'h16ba: color = 2'b10;
      13'h16bb: color = 2'b10;
      13'h16bc: color = 2'b10;
      13'h16bd: color = 2'b10;
      13'h16be: color = 2'b10;
      13'h16bf: color = 2'b10;
      13'h16c0: color = 2'b10;
      13'h16c1: color = 2'b10;
      13'h16c2: color = 2'b10;
      13'h16c3: color = 2'b10;
      13'h16c4: color = 2'b10;
      13'h16c5: color = 2'b10;
      13'h16c6: color = 2'b10;
      13'h16c7: color = 2'b10;
      13'h16c8: color = 2'b10;
      13'h16c9: color = 2'b10;
      13'h16ca: color = 2'b10;
      13'h16cb: color = 2'b10;
      13'h16cc: color = 2'b10;
      13'h16cd: color = 2'b10;
      13'h16ce: color = 2'b10;
      13'h16cf: color = 2'b10;
      13'h16d0: color = 2'b10;
      13'h16d1: color = 2'b10;
      13'h16d2: color = 2'b10;
      13'h16d3: color = 2'b10;
      13'h16d4: color = 2'b10;
      13'h16d5: color = 2'b10;
      13'h16d6: color = 2'b10;
      13'h16d7: color = 2'b10;
      13'h16d8: color = 2'b10;
      13'h16d9: color = 2'b10;
      13'h16da: color = 2'b10;
      13'h16db: color = 2'b10;
      13'h16dc: color = 2'b01;
      13'h16dd: color = 2'b01;
      13'h16de: color = 2'b00;
      13'h16df: color = 2'b00;
      13'h16e0: color = 2'b11;
      13'h16e1: color = 2'b11;
      13'h16e2: color = 2'b11;
      13'h16e3: color = 2'b11;
      13'h16e4: color = 2'b00;
      13'h16e5: color = 2'b00;
      13'h16e6: color = 2'b11;
      13'h16e7: color = 2'b11;
      13'h16e8: color = 2'b11;
      13'h16e9: color = 2'b11;
      13'h16ea: color = 2'b11;
      13'h16eb: color = 2'b11;
      13'h16ec: color = 2'b11;
      13'h16ed: color = 2'b11;
      13'h16ee: color = 2'b11;
      13'h16ef: color = 2'b11;
      13'h16f0: color = 2'b11;
      13'h16f1: color = 2'b11;
      13'h16f2: color = 2'b11;
      13'h16f3: color = 2'b11;
      13'h16f4: color = 2'b11;
      13'h16f5: color = 2'b11;
      13'h16f6: color = 2'b11;
      13'h16f7: color = 2'b11;
      13'h16f8: color = 2'b11;
      13'h16f9: color = 2'b11;
      13'h16fa: color = 2'b00;
      13'h16fb: color = 2'b00;
      13'h16fc: color = 2'b11;
      13'h16fd: color = 2'b11;
      13'h16fe: color = 2'b11;
      13'h16ff: color = 2'b11;
      13'h1700: color = 2'b11;
      13'h1701: color = 2'b11;
      13'h1702: color = 2'b11;
      13'h1703: color = 2'b11;
      13'h1704: color = 2'b00;
      13'h1705: color = 2'b00;
      13'h1706: color = 2'b11;
      13'h1707: color = 2'b11;
      13'h1708: color = 2'b11;
      13'h1709: color = 2'b11;
      13'h170a: color = 2'b10;
      13'h170b: color = 2'b10;
      13'h170c: color = 2'b10;
      13'h170d: color = 2'b10;
      13'h170e: color = 2'b10;
      13'h170f: color = 2'b10;
      13'h1710: color = 2'b10;
      13'h1711: color = 2'b10;
      13'h1712: color = 2'b10;
      13'h1713: color = 2'b10;
      13'h1714: color = 2'b10;
      13'h1715: color = 2'b10;
      13'h1716: color = 2'b11;
      13'h1717: color = 2'b11;
      13'h1718: color = 2'b11;
      13'h1719: color = 2'b11;
      13'h171a: color = 2'b00;
      13'h171b: color = 2'b00;
      13'h171c: color = 2'b11;
      13'h171d: color = 2'b11;
      13'h171e: color = 2'b11;
      13'h171f: color = 2'b11;
      13'h1720: color = 2'b00;
      13'h1721: color = 2'b00;
      13'h1722: color = 2'b00;
      13'h1723: color = 2'b00;
      13'h1724: color = 2'b01;
      13'h1725: color = 2'b01;
      13'h1726: color = 2'b01;
      13'h1727: color = 2'b01;
      13'h1728: color = 2'b01;
      13'h1729: color = 2'b01;
      13'h172a: color = 2'b01;
      13'h172b: color = 2'b01;
      13'h172c: color = 2'b01;
      13'h172d: color = 2'b01;
      13'h172e: color = 2'b01;
      13'h172f: color = 2'b01;
      13'h1730: color = 2'b01;
      13'h1731: color = 2'b01;
      13'h1732: color = 2'b01;
      13'h1733: color = 2'b01;
      13'h1734: color = 2'b01;
      13'h1735: color = 2'b01;
      13'h1736: color = 2'b01;
      13'h1737: color = 2'b01;
      13'h1738: color = 2'b01;
      13'h1739: color = 2'b01;
      13'h173a: color = 2'b01;
      13'h173b: color = 2'b01;
      13'h173c: color = 2'b01;
      13'h173d: color = 2'b01;
      13'h173e: color = 2'b01;
      13'h173f: color = 2'b01;
      13'h1740: color = 2'b01;
      13'h1741: color = 2'b01;
      13'h1742: color = 2'b01;
      13'h1743: color = 2'b01;
      13'h1744: color = 2'b01;
      13'h1745: color = 2'b01;
      13'h1746: color = 2'b01;
      13'h1747: color = 2'b01;
      13'h1748: color = 2'b01;
      13'h1749: color = 2'b01;
      13'h174a: color = 2'b01;
      13'h174b: color = 2'b01;
      13'h174c: color = 2'b01;
      13'h174d: color = 2'b01;
      13'h174e: color = 2'b01;
      13'h174f: color = 2'b01;
      13'h1750: color = 2'b01;
      13'h1751: color = 2'b01;
      13'h1752: color = 2'b01;
      13'h1753: color = 2'b01;
      13'h1754: color = 2'b01;
      13'h1755: color = 2'b01;
      13'h1756: color = 2'b01;
      13'h1757: color = 2'b01;
      13'h1758: color = 2'b01;
      13'h1759: color = 2'b01;
      13'h175a: color = 2'b01;
      13'h175b: color = 2'b01;
      13'h175c: color = 2'b00;
      13'h175d: color = 2'b00;
      13'h175e: color = 2'b00;
      13'h175f: color = 2'b00;
      13'h1760: color = 2'b11;
      13'h1761: color = 2'b11;
      13'h1762: color = 2'b11;
      13'h1763: color = 2'b11;
      13'h1764: color = 2'b00;
      13'h1765: color = 2'b00;
      13'h1766: color = 2'b11;
      13'h1767: color = 2'b11;
      13'h1768: color = 2'b11;
      13'h1769: color = 2'b11;
      13'h176a: color = 2'b10;
      13'h176b: color = 2'b10;
      13'h176c: color = 2'b10;
      13'h176d: color = 2'b10;
      13'h176e: color = 2'b10;
      13'h176f: color = 2'b10;
      13'h1770: color = 2'b10;
      13'h1771: color = 2'b10;
      13'h1772: color = 2'b10;
      13'h1773: color = 2'b10;
      13'h1774: color = 2'b10;
      13'h1775: color = 2'b10;
      13'h1776: color = 2'b11;
      13'h1777: color = 2'b11;
      13'h1778: color = 2'b11;
      13'h1779: color = 2'b11;
      13'h177a: color = 2'b00;
      13'h177b: color = 2'b00;
      13'h177c: color = 2'b11;
      13'h177d: color = 2'b11;
      13'h177e: color = 2'b11;
      13'h177f: color = 2'b11;
      13'h1780: color = 2'b11;
      13'h1781: color = 2'b11;
      13'h1782: color = 2'b11;
      13'h1783: color = 2'b11;
      13'h1784: color = 2'b00;
      13'h1785: color = 2'b00;
      13'h1786: color = 2'b11;
      13'h1787: color = 2'b11;
      13'h1788: color = 2'b11;
      13'h1789: color = 2'b11;
      13'h178a: color = 2'b10;
      13'h178b: color = 2'b10;
      13'h178c: color = 2'b10;
      13'h178d: color = 2'b10;
      13'h178e: color = 2'b10;
      13'h178f: color = 2'b10;
      13'h1790: color = 2'b10;
      13'h1791: color = 2'b10;
      13'h1792: color = 2'b10;
      13'h1793: color = 2'b10;
      13'h1794: color = 2'b10;
      13'h1795: color = 2'b10;
      13'h1796: color = 2'b11;
      13'h1797: color = 2'b11;
      13'h1798: color = 2'b11;
      13'h1799: color = 2'b11;
      13'h179a: color = 2'b00;
      13'h179b: color = 2'b00;
      13'h179c: color = 2'b11;
      13'h179d: color = 2'b11;
      13'h179e: color = 2'b11;
      13'h179f: color = 2'b11;
      13'h17a0: color = 2'b00;
      13'h17a1: color = 2'b00;
      13'h17a2: color = 2'b00;
      13'h17a3: color = 2'b00;
      13'h17a4: color = 2'b01;
      13'h17a5: color = 2'b01;
      13'h17a6: color = 2'b01;
      13'h17a7: color = 2'b01;
      13'h17a8: color = 2'b01;
      13'h17a9: color = 2'b01;
      13'h17aa: color = 2'b01;
      13'h17ab: color = 2'b01;
      13'h17ac: color = 2'b01;
      13'h17ad: color = 2'b01;
      13'h17ae: color = 2'b01;
      13'h17af: color = 2'b01;
      13'h17b0: color = 2'b01;
      13'h17b1: color = 2'b01;
      13'h17b2: color = 2'b01;
      13'h17b3: color = 2'b01;
      13'h17b4: color = 2'b01;
      13'h17b5: color = 2'b01;
      13'h17b6: color = 2'b01;
      13'h17b7: color = 2'b01;
      13'h17b8: color = 2'b01;
      13'h17b9: color = 2'b01;
      13'h17ba: color = 2'b01;
      13'h17bb: color = 2'b01;
      13'h17bc: color = 2'b01;
      13'h17bd: color = 2'b01;
      13'h17be: color = 2'b01;
      13'h17bf: color = 2'b01;
      13'h17c0: color = 2'b01;
      13'h17c1: color = 2'b01;
      13'h17c2: color = 2'b01;
      13'h17c3: color = 2'b01;
      13'h17c4: color = 2'b01;
      13'h17c5: color = 2'b01;
      13'h17c6: color = 2'b01;
      13'h17c7: color = 2'b01;
      13'h17c8: color = 2'b01;
      13'h17c9: color = 2'b01;
      13'h17ca: color = 2'b01;
      13'h17cb: color = 2'b01;
      13'h17cc: color = 2'b01;
      13'h17cd: color = 2'b01;
      13'h17ce: color = 2'b01;
      13'h17cf: color = 2'b01;
      13'h17d0: color = 2'b01;
      13'h17d1: color = 2'b01;
      13'h17d2: color = 2'b01;
      13'h17d3: color = 2'b01;
      13'h17d4: color = 2'b01;
      13'h17d5: color = 2'b01;
      13'h17d6: color = 2'b01;
      13'h17d7: color = 2'b01;
      13'h17d8: color = 2'b01;
      13'h17d9: color = 2'b01;
      13'h17da: color = 2'b01;
      13'h17db: color = 2'b01;
      13'h17dc: color = 2'b00;
      13'h17dd: color = 2'b00;
      13'h17de: color = 2'b00;
      13'h17df: color = 2'b00;
      13'h17e0: color = 2'b11;
      13'h17e1: color = 2'b11;
      13'h17e2: color = 2'b11;
      13'h17e3: color = 2'b11;
      13'h17e4: color = 2'b00;
      13'h17e5: color = 2'b00;
      13'h17e6: color = 2'b11;
      13'h17e7: color = 2'b11;
      13'h17e8: color = 2'b11;
      13'h17e9: color = 2'b11;
      13'h17ea: color = 2'b10;
      13'h17eb: color = 2'b10;
      13'h17ec: color = 2'b10;
      13'h17ed: color = 2'b10;
      13'h17ee: color = 2'b10;
      13'h17ef: color = 2'b10;
      13'h17f0: color = 2'b10;
      13'h17f1: color = 2'b10;
      13'h17f2: color = 2'b10;
      13'h17f3: color = 2'b10;
      13'h17f4: color = 2'b10;
      13'h17f5: color = 2'b10;
      13'h17f6: color = 2'b11;
      13'h17f7: color = 2'b11;
      13'h17f8: color = 2'b11;
      13'h17f9: color = 2'b11;
      13'h17fa: color = 2'b00;
      13'h17fb: color = 2'b00;
      13'h17fc: color = 2'b11;
      13'h17fd: color = 2'b11;
      13'h17fe: color = 2'b11;
      13'h17ff: color = 2'b11;
      13'h1800: color = 2'b11;
      13'h1801: color = 2'b11;
      13'h1802: color = 2'b11;
      13'h1803: color = 2'b11;
      13'h1804: color = 2'b00;
      13'h1805: color = 2'b00;
      13'h1806: color = 2'b11;
      13'h1807: color = 2'b11;
      13'h1808: color = 2'b11;
      13'h1809: color = 2'b11;
      13'h180a: color = 2'b10;
      13'h180b: color = 2'b10;
      13'h180c: color = 2'b10;
      13'h180d: color = 2'b10;
      13'h180e: color = 2'b10;
      13'h180f: color = 2'b10;
      13'h1810: color = 2'b10;
      13'h1811: color = 2'b10;
      13'h1812: color = 2'b10;
      13'h1813: color = 2'b10;
      13'h1814: color = 2'b10;
      13'h1815: color = 2'b10;
      13'h1816: color = 2'b11;
      13'h1817: color = 2'b11;
      13'h1818: color = 2'b11;
      13'h1819: color = 2'b11;
      13'h181a: color = 2'b00;
      13'h181b: color = 2'b00;
      13'h181c: color = 2'b11;
      13'h181d: color = 2'b11;
      13'h181e: color = 2'b11;
      13'h181f: color = 2'b11;
      13'h1820: color = 2'b00;
      13'h1821: color = 2'b00;
      13'h1822: color = 2'b00;
      13'h1823: color = 2'b00;
      13'h1824: color = 2'b00;
      13'h1825: color = 2'b00;
      13'h1826: color = 2'b00;
      13'h1827: color = 2'b00;
      13'h1828: color = 2'b00;
      13'h1829: color = 2'b00;
      13'h182a: color = 2'b00;
      13'h182b: color = 2'b00;
      13'h182c: color = 2'b00;
      13'h182d: color = 2'b00;
      13'h182e: color = 2'b00;
      13'h182f: color = 2'b00;
      13'h1830: color = 2'b00;
      13'h1831: color = 2'b00;
      13'h1832: color = 2'b00;
      13'h1833: color = 2'b00;
      13'h1834: color = 2'b00;
      13'h1835: color = 2'b00;
      13'h1836: color = 2'b00;
      13'h1837: color = 2'b00;
      13'h1838: color = 2'b00;
      13'h1839: color = 2'b00;
      13'h183a: color = 2'b00;
      13'h183b: color = 2'b00;
      13'h183c: color = 2'b00;
      13'h183d: color = 2'b00;
      13'h183e: color = 2'b00;
      13'h183f: color = 2'b00;
      13'h1840: color = 2'b00;
      13'h1841: color = 2'b00;
      13'h1842: color = 2'b00;
      13'h1843: color = 2'b00;
      13'h1844: color = 2'b00;
      13'h1845: color = 2'b00;
      13'h1846: color = 2'b00;
      13'h1847: color = 2'b00;
      13'h1848: color = 2'b00;
      13'h1849: color = 2'b00;
      13'h184a: color = 2'b00;
      13'h184b: color = 2'b00;
      13'h184c: color = 2'b00;
      13'h184d: color = 2'b00;
      13'h184e: color = 2'b00;
      13'h184f: color = 2'b00;
      13'h1850: color = 2'b00;
      13'h1851: color = 2'b00;
      13'h1852: color = 2'b00;
      13'h1853: color = 2'b00;
      13'h1854: color = 2'b00;
      13'h1855: color = 2'b00;
      13'h1856: color = 2'b00;
      13'h1857: color = 2'b00;
      13'h1858: color = 2'b00;
      13'h1859: color = 2'b00;
      13'h185a: color = 2'b00;
      13'h185b: color = 2'b00;
      13'h185c: color = 2'b00;
      13'h185d: color = 2'b00;
      13'h185e: color = 2'b00;
      13'h185f: color = 2'b00;
      13'h1860: color = 2'b11;
      13'h1861: color = 2'b11;
      13'h1862: color = 2'b11;
      13'h1863: color = 2'b11;
      13'h1864: color = 2'b00;
      13'h1865: color = 2'b00;
      13'h1866: color = 2'b11;
      13'h1867: color = 2'b11;
      13'h1868: color = 2'b11;
      13'h1869: color = 2'b11;
      13'h186a: color = 2'b10;
      13'h186b: color = 2'b10;
      13'h186c: color = 2'b10;
      13'h186d: color = 2'b10;
      13'h186e: color = 2'b10;
      13'h186f: color = 2'b10;
      13'h1870: color = 2'b10;
      13'h1871: color = 2'b10;
      13'h1872: color = 2'b10;
      13'h1873: color = 2'b10;
      13'h1874: color = 2'b10;
      13'h1875: color = 2'b10;
      13'h1876: color = 2'b11;
      13'h1877: color = 2'b11;
      13'h1878: color = 2'b11;
      13'h1879: color = 2'b11;
      13'h187a: color = 2'b00;
      13'h187b: color = 2'b00;
      13'h187c: color = 2'b11;
      13'h187d: color = 2'b11;
      13'h187e: color = 2'b11;
      13'h187f: color = 2'b11;
      13'h1880: color = 2'b11;
      13'h1881: color = 2'b11;
      13'h1882: color = 2'b11;
      13'h1883: color = 2'b11;
      13'h1884: color = 2'b00;
      13'h1885: color = 2'b00;
      13'h1886: color = 2'b11;
      13'h1887: color = 2'b11;
      13'h1888: color = 2'b11;
      13'h1889: color = 2'b11;
      13'h188a: color = 2'b10;
      13'h188b: color = 2'b10;
      13'h188c: color = 2'b10;
      13'h188d: color = 2'b10;
      13'h188e: color = 2'b10;
      13'h188f: color = 2'b10;
      13'h1890: color = 2'b10;
      13'h1891: color = 2'b10;
      13'h1892: color = 2'b10;
      13'h1893: color = 2'b10;
      13'h1894: color = 2'b10;
      13'h1895: color = 2'b10;
      13'h1896: color = 2'b11;
      13'h1897: color = 2'b11;
      13'h1898: color = 2'b11;
      13'h1899: color = 2'b11;
      13'h189a: color = 2'b00;
      13'h189b: color = 2'b00;
      13'h189c: color = 2'b11;
      13'h189d: color = 2'b11;
      13'h189e: color = 2'b11;
      13'h189f: color = 2'b11;
      13'h18a0: color = 2'b00;
      13'h18a1: color = 2'b00;
      13'h18a2: color = 2'b00;
      13'h18a3: color = 2'b00;
      13'h18a4: color = 2'b00;
      13'h18a5: color = 2'b00;
      13'h18a6: color = 2'b00;
      13'h18a7: color = 2'b00;
      13'h18a8: color = 2'b00;
      13'h18a9: color = 2'b00;
      13'h18aa: color = 2'b00;
      13'h18ab: color = 2'b00;
      13'h18ac: color = 2'b00;
      13'h18ad: color = 2'b00;
      13'h18ae: color = 2'b00;
      13'h18af: color = 2'b00;
      13'h18b0: color = 2'b00;
      13'h18b1: color = 2'b00;
      13'h18b2: color = 2'b00;
      13'h18b3: color = 2'b00;
      13'h18b4: color = 2'b00;
      13'h18b5: color = 2'b00;
      13'h18b6: color = 2'b00;
      13'h18b7: color = 2'b00;
      13'h18b8: color = 2'b00;
      13'h18b9: color = 2'b00;
      13'h18ba: color = 2'b00;
      13'h18bb: color = 2'b00;
      13'h18bc: color = 2'b00;
      13'h18bd: color = 2'b00;
      13'h18be: color = 2'b00;
      13'h18bf: color = 2'b00;
      13'h18c0: color = 2'b00;
      13'h18c1: color = 2'b00;
      13'h18c2: color = 2'b00;
      13'h18c3: color = 2'b00;
      13'h18c4: color = 2'b00;
      13'h18c5: color = 2'b00;
      13'h18c6: color = 2'b00;
      13'h18c7: color = 2'b00;
      13'h18c8: color = 2'b00;
      13'h18c9: color = 2'b00;
      13'h18ca: color = 2'b00;
      13'h18cb: color = 2'b00;
      13'h18cc: color = 2'b00;
      13'h18cd: color = 2'b00;
      13'h18ce: color = 2'b00;
      13'h18cf: color = 2'b00;
      13'h18d0: color = 2'b00;
      13'h18d1: color = 2'b00;
      13'h18d2: color = 2'b00;
      13'h18d3: color = 2'b00;
      13'h18d4: color = 2'b00;
      13'h18d5: color = 2'b00;
      13'h18d6: color = 2'b00;
      13'h18d7: color = 2'b00;
      13'h18d8: color = 2'b00;
      13'h18d9: color = 2'b00;
      13'h18da: color = 2'b00;
      13'h18db: color = 2'b00;
      13'h18dc: color = 2'b00;
      13'h18dd: color = 2'b00;
      13'h18de: color = 2'b00;
      13'h18df: color = 2'b00;
      13'h18e0: color = 2'b11;
      13'h18e1: color = 2'b11;
      13'h18e2: color = 2'b11;
      13'h18e3: color = 2'b11;
      13'h18e4: color = 2'b00;
      13'h18e5: color = 2'b00;
      13'h18e6: color = 2'b11;
      13'h18e7: color = 2'b11;
      13'h18e8: color = 2'b11;
      13'h18e9: color = 2'b11;
      13'h18ea: color = 2'b10;
      13'h18eb: color = 2'b10;
      13'h18ec: color = 2'b10;
      13'h18ed: color = 2'b10;
      13'h18ee: color = 2'b10;
      13'h18ef: color = 2'b10;
      13'h18f0: color = 2'b10;
      13'h18f1: color = 2'b10;
      13'h18f2: color = 2'b10;
      13'h18f3: color = 2'b10;
      13'h18f4: color = 2'b10;
      13'h18f5: color = 2'b10;
      13'h18f6: color = 2'b11;
      13'h18f7: color = 2'b11;
      13'h18f8: color = 2'b11;
      13'h18f9: color = 2'b11;
      13'h18fa: color = 2'b00;
      13'h18fb: color = 2'b00;
      13'h18fc: color = 2'b11;
      13'h18fd: color = 2'b11;
      13'h18fe: color = 2'b11;
      13'h18ff: color = 2'b11;
      13'h1900: color = 2'b11;
      13'h1901: color = 2'b11;
      13'h1902: color = 2'b10;
      13'h1903: color = 2'b10;
      13'h1904: color = 2'b00;
      13'h1905: color = 2'b00;
      13'h1906: color = 2'b11;
      13'h1907: color = 2'b11;
      13'h1908: color = 2'b11;
      13'h1909: color = 2'b11;
      13'h190a: color = 2'b10;
      13'h190b: color = 2'b10;
      13'h190c: color = 2'b10;
      13'h190d: color = 2'b10;
      13'h190e: color = 2'b10;
      13'h190f: color = 2'b10;
      13'h1910: color = 2'b10;
      13'h1911: color = 2'b10;
      13'h1912: color = 2'b10;
      13'h1913: color = 2'b10;
      13'h1914: color = 2'b10;
      13'h1915: color = 2'b10;
      13'h1916: color = 2'b11;
      13'h1917: color = 2'b11;
      13'h1918: color = 2'b11;
      13'h1919: color = 2'b11;
      13'h191a: color = 2'b00;
      13'h191b: color = 2'b00;
      13'h191c: color = 2'b11;
      13'h191d: color = 2'b11;
      13'h191e: color = 2'b11;
      13'h191f: color = 2'b11;
      13'h1920: color = 2'b00;
      13'h1921: color = 2'b00;
      13'h1922: color = 2'b01;
      13'h1923: color = 2'b01;
      13'h1924: color = 2'b01;
      13'h1925: color = 2'b01;
      13'h1926: color = 2'b01;
      13'h1927: color = 2'b01;
      13'h1928: color = 2'b01;
      13'h1929: color = 2'b01;
      13'h192a: color = 2'b01;
      13'h192b: color = 2'b01;
      13'h192c: color = 2'b01;
      13'h192d: color = 2'b01;
      13'h192e: color = 2'b01;
      13'h192f: color = 2'b01;
      13'h1930: color = 2'b01;
      13'h1931: color = 2'b01;
      13'h1932: color = 2'b01;
      13'h1933: color = 2'b01;
      13'h1934: color = 2'b01;
      13'h1935: color = 2'b01;
      13'h1936: color = 2'b01;
      13'h1937: color = 2'b01;
      13'h1938: color = 2'b01;
      13'h1939: color = 2'b01;
      13'h193a: color = 2'b01;
      13'h193b: color = 2'b01;
      13'h193c: color = 2'b01;
      13'h193d: color = 2'b01;
      13'h193e: color = 2'b01;
      13'h193f: color = 2'b01;
      13'h1940: color = 2'b01;
      13'h1941: color = 2'b01;
      13'h1942: color = 2'b01;
      13'h1943: color = 2'b01;
      13'h1944: color = 2'b01;
      13'h1945: color = 2'b01;
      13'h1946: color = 2'b01;
      13'h1947: color = 2'b01;
      13'h1948: color = 2'b01;
      13'h1949: color = 2'b01;
      13'h194a: color = 2'b01;
      13'h194b: color = 2'b01;
      13'h194c: color = 2'b01;
      13'h194d: color = 2'b01;
      13'h194e: color = 2'b01;
      13'h194f: color = 2'b01;
      13'h1950: color = 2'b01;
      13'h1951: color = 2'b01;
      13'h1952: color = 2'b01;
      13'h1953: color = 2'b01;
      13'h1954: color = 2'b01;
      13'h1955: color = 2'b01;
      13'h1956: color = 2'b01;
      13'h1957: color = 2'b01;
      13'h1958: color = 2'b01;
      13'h1959: color = 2'b01;
      13'h195a: color = 2'b01;
      13'h195b: color = 2'b01;
      13'h195c: color = 2'b01;
      13'h195d: color = 2'b01;
      13'h195e: color = 2'b00;
      13'h195f: color = 2'b00;
      13'h1960: color = 2'b11;
      13'h1961: color = 2'b11;
      13'h1962: color = 2'b10;
      13'h1963: color = 2'b10;
      13'h1964: color = 2'b00;
      13'h1965: color = 2'b00;
      13'h1966: color = 2'b11;
      13'h1967: color = 2'b11;
      13'h1968: color = 2'b11;
      13'h1969: color = 2'b11;
      13'h196a: color = 2'b10;
      13'h196b: color = 2'b10;
      13'h196c: color = 2'b10;
      13'h196d: color = 2'b10;
      13'h196e: color = 2'b10;
      13'h196f: color = 2'b10;
      13'h1970: color = 2'b10;
      13'h1971: color = 2'b10;
      13'h1972: color = 2'b10;
      13'h1973: color = 2'b10;
      13'h1974: color = 2'b10;
      13'h1975: color = 2'b10;
      13'h1976: color = 2'b11;
      13'h1977: color = 2'b11;
      13'h1978: color = 2'b11;
      13'h1979: color = 2'b11;
      13'h197a: color = 2'b00;
      13'h197b: color = 2'b00;
      13'h197c: color = 2'b11;
      13'h197d: color = 2'b11;
      13'h197e: color = 2'b11;
      13'h197f: color = 2'b11;
      13'h1980: color = 2'b11;
      13'h1981: color = 2'b11;
      13'h1982: color = 2'b10;
      13'h1983: color = 2'b10;
      13'h1984: color = 2'b00;
      13'h1985: color = 2'b00;
      13'h1986: color = 2'b11;
      13'h1987: color = 2'b11;
      13'h1988: color = 2'b11;
      13'h1989: color = 2'b11;
      13'h198a: color = 2'b10;
      13'h198b: color = 2'b10;
      13'h198c: color = 2'b10;
      13'h198d: color = 2'b10;
      13'h198e: color = 2'b10;
      13'h198f: color = 2'b10;
      13'h1990: color = 2'b10;
      13'h1991: color = 2'b10;
      13'h1992: color = 2'b10;
      13'h1993: color = 2'b10;
      13'h1994: color = 2'b10;
      13'h1995: color = 2'b10;
      13'h1996: color = 2'b11;
      13'h1997: color = 2'b11;
      13'h1998: color = 2'b11;
      13'h1999: color = 2'b11;
      13'h199a: color = 2'b00;
      13'h199b: color = 2'b00;
      13'h199c: color = 2'b11;
      13'h199d: color = 2'b11;
      13'h199e: color = 2'b11;
      13'h199f: color = 2'b11;
      13'h19a0: color = 2'b00;
      13'h19a1: color = 2'b00;
      13'h19a2: color = 2'b01;
      13'h19a3: color = 2'b01;
      13'h19a4: color = 2'b01;
      13'h19a5: color = 2'b01;
      13'h19a6: color = 2'b01;
      13'h19a7: color = 2'b01;
      13'h19a8: color = 2'b01;
      13'h19a9: color = 2'b01;
      13'h19aa: color = 2'b01;
      13'h19ab: color = 2'b01;
      13'h19ac: color = 2'b01;
      13'h19ad: color = 2'b01;
      13'h19ae: color = 2'b01;
      13'h19af: color = 2'b01;
      13'h19b0: color = 2'b01;
      13'h19b1: color = 2'b01;
      13'h19b2: color = 2'b01;
      13'h19b3: color = 2'b01;
      13'h19b4: color = 2'b01;
      13'h19b5: color = 2'b01;
      13'h19b6: color = 2'b01;
      13'h19b7: color = 2'b01;
      13'h19b8: color = 2'b01;
      13'h19b9: color = 2'b01;
      13'h19ba: color = 2'b01;
      13'h19bb: color = 2'b01;
      13'h19bc: color = 2'b01;
      13'h19bd: color = 2'b01;
      13'h19be: color = 2'b01;
      13'h19bf: color = 2'b01;
      13'h19c0: color = 2'b01;
      13'h19c1: color = 2'b01;
      13'h19c2: color = 2'b01;
      13'h19c3: color = 2'b01;
      13'h19c4: color = 2'b01;
      13'h19c5: color = 2'b01;
      13'h19c6: color = 2'b01;
      13'h19c7: color = 2'b01;
      13'h19c8: color = 2'b01;
      13'h19c9: color = 2'b01;
      13'h19ca: color = 2'b01;
      13'h19cb: color = 2'b01;
      13'h19cc: color = 2'b01;
      13'h19cd: color = 2'b01;
      13'h19ce: color = 2'b01;
      13'h19cf: color = 2'b01;
      13'h19d0: color = 2'b01;
      13'h19d1: color = 2'b01;
      13'h19d2: color = 2'b01;
      13'h19d3: color = 2'b01;
      13'h19d4: color = 2'b01;
      13'h19d5: color = 2'b01;
      13'h19d6: color = 2'b01;
      13'h19d7: color = 2'b01;
      13'h19d8: color = 2'b01;
      13'h19d9: color = 2'b01;
      13'h19da: color = 2'b01;
      13'h19db: color = 2'b01;
      13'h19dc: color = 2'b01;
      13'h19dd: color = 2'b01;
      13'h19de: color = 2'b00;
      13'h19df: color = 2'b00;
      13'h19e0: color = 2'b11;
      13'h19e1: color = 2'b11;
      13'h19e2: color = 2'b10;
      13'h19e3: color = 2'b10;
      13'h19e4: color = 2'b00;
      13'h19e5: color = 2'b00;
      13'h19e6: color = 2'b11;
      13'h19e7: color = 2'b11;
      13'h19e8: color = 2'b11;
      13'h19e9: color = 2'b11;
      13'h19ea: color = 2'b10;
      13'h19eb: color = 2'b10;
      13'h19ec: color = 2'b10;
      13'h19ed: color = 2'b10;
      13'h19ee: color = 2'b10;
      13'h19ef: color = 2'b10;
      13'h19f0: color = 2'b10;
      13'h19f1: color = 2'b10;
      13'h19f2: color = 2'b10;
      13'h19f3: color = 2'b10;
      13'h19f4: color = 2'b10;
      13'h19f5: color = 2'b10;
      13'h19f6: color = 2'b11;
      13'h19f7: color = 2'b11;
      13'h19f8: color = 2'b11;
      13'h19f9: color = 2'b11;
      13'h19fa: color = 2'b00;
      13'h19fb: color = 2'b00;
      13'h19fc: color = 2'b11;
      13'h19fd: color = 2'b11;
      13'h19fe: color = 2'b11;
      13'h19ff: color = 2'b11;
      13'h1a00: color = 2'b10;
      13'h1a01: color = 2'b10;
      13'h1a02: color = 2'b11;
      13'h1a03: color = 2'b11;
      13'h1a04: color = 2'b00;
      13'h1a05: color = 2'b00;
      13'h1a06: color = 2'b11;
      13'h1a07: color = 2'b11;
      13'h1a08: color = 2'b11;
      13'h1a09: color = 2'b11;
      13'h1a0a: color = 2'b11;
      13'h1a0b: color = 2'b11;
      13'h1a0c: color = 2'b11;
      13'h1a0d: color = 2'b11;
      13'h1a0e: color = 2'b11;
      13'h1a0f: color = 2'b11;
      13'h1a10: color = 2'b11;
      13'h1a11: color = 2'b11;
      13'h1a12: color = 2'b11;
      13'h1a13: color = 2'b11;
      13'h1a14: color = 2'b11;
      13'h1a15: color = 2'b11;
      13'h1a16: color = 2'b11;
      13'h1a17: color = 2'b11;
      13'h1a18: color = 2'b11;
      13'h1a19: color = 2'b11;
      13'h1a1a: color = 2'b00;
      13'h1a1b: color = 2'b00;
      13'h1a1c: color = 2'b10;
      13'h1a1d: color = 2'b10;
      13'h1a1e: color = 2'b11;
      13'h1a1f: color = 2'b11;
      13'h1a20: color = 2'b10;
      13'h1a21: color = 2'b10;
      13'h1a22: color = 2'b00;
      13'h1a23: color = 2'b00;
      13'h1a24: color = 2'b00;
      13'h1a25: color = 2'b00;
      13'h1a26: color = 2'b00;
      13'h1a27: color = 2'b00;
      13'h1a28: color = 2'b00;
      13'h1a29: color = 2'b00;
      13'h1a2a: color = 2'b00;
      13'h1a2b: color = 2'b00;
      13'h1a2c: color = 2'b00;
      13'h1a2d: color = 2'b00;
      13'h1a2e: color = 2'b00;
      13'h1a2f: color = 2'b00;
      13'h1a30: color = 2'b00;
      13'h1a31: color = 2'b00;
      13'h1a32: color = 2'b00;
      13'h1a33: color = 2'b00;
      13'h1a34: color = 2'b00;
      13'h1a35: color = 2'b00;
      13'h1a36: color = 2'b00;
      13'h1a37: color = 2'b00;
      13'h1a38: color = 2'b00;
      13'h1a39: color = 2'b00;
      13'h1a3a: color = 2'b00;
      13'h1a3b: color = 2'b00;
      13'h1a3c: color = 2'b00;
      13'h1a3d: color = 2'b00;
      13'h1a3e: color = 2'b00;
      13'h1a3f: color = 2'b00;
      13'h1a40: color = 2'b00;
      13'h1a41: color = 2'b00;
      13'h1a42: color = 2'b00;
      13'h1a43: color = 2'b00;
      13'h1a44: color = 2'b00;
      13'h1a45: color = 2'b00;
      13'h1a46: color = 2'b00;
      13'h1a47: color = 2'b00;
      13'h1a48: color = 2'b00;
      13'h1a49: color = 2'b00;
      13'h1a4a: color = 2'b00;
      13'h1a4b: color = 2'b00;
      13'h1a4c: color = 2'b00;
      13'h1a4d: color = 2'b00;
      13'h1a4e: color = 2'b00;
      13'h1a4f: color = 2'b00;
      13'h1a50: color = 2'b00;
      13'h1a51: color = 2'b00;
      13'h1a52: color = 2'b00;
      13'h1a53: color = 2'b00;
      13'h1a54: color = 2'b00;
      13'h1a55: color = 2'b00;
      13'h1a56: color = 2'b00;
      13'h1a57: color = 2'b00;
      13'h1a58: color = 2'b00;
      13'h1a59: color = 2'b00;
      13'h1a5a: color = 2'b00;
      13'h1a5b: color = 2'b00;
      13'h1a5c: color = 2'b00;
      13'h1a5d: color = 2'b00;
      13'h1a5e: color = 2'b11;
      13'h1a5f: color = 2'b11;
      13'h1a60: color = 2'b10;
      13'h1a61: color = 2'b10;
      13'h1a62: color = 2'b11;
      13'h1a63: color = 2'b11;
      13'h1a64: color = 2'b00;
      13'h1a65: color = 2'b00;
      13'h1a66: color = 2'b11;
      13'h1a67: color = 2'b11;
      13'h1a68: color = 2'b11;
      13'h1a69: color = 2'b11;
      13'h1a6a: color = 2'b11;
      13'h1a6b: color = 2'b11;
      13'h1a6c: color = 2'b11;
      13'h1a6d: color = 2'b11;
      13'h1a6e: color = 2'b11;
      13'h1a6f: color = 2'b11;
      13'h1a70: color = 2'b11;
      13'h1a71: color = 2'b11;
      13'h1a72: color = 2'b11;
      13'h1a73: color = 2'b11;
      13'h1a74: color = 2'b11;
      13'h1a75: color = 2'b11;
      13'h1a76: color = 2'b11;
      13'h1a77: color = 2'b11;
      13'h1a78: color = 2'b11;
      13'h1a79: color = 2'b11;
      13'h1a7a: color = 2'b00;
      13'h1a7b: color = 2'b00;
      13'h1a7c: color = 2'b10;
      13'h1a7d: color = 2'b10;
      13'h1a7e: color = 2'b11;
      13'h1a7f: color = 2'b11;
      13'h1a80: color = 2'b10;
      13'h1a81: color = 2'b10;
      13'h1a82: color = 2'b11;
      13'h1a83: color = 2'b11;
      13'h1a84: color = 2'b00;
      13'h1a85: color = 2'b00;
      13'h1a86: color = 2'b11;
      13'h1a87: color = 2'b11;
      13'h1a88: color = 2'b11;
      13'h1a89: color = 2'b11;
      13'h1a8a: color = 2'b11;
      13'h1a8b: color = 2'b11;
      13'h1a8c: color = 2'b11;
      13'h1a8d: color = 2'b11;
      13'h1a8e: color = 2'b11;
      13'h1a8f: color = 2'b11;
      13'h1a90: color = 2'b11;
      13'h1a91: color = 2'b11;
      13'h1a92: color = 2'b11;
      13'h1a93: color = 2'b11;
      13'h1a94: color = 2'b11;
      13'h1a95: color = 2'b11;
      13'h1a96: color = 2'b11;
      13'h1a97: color = 2'b11;
      13'h1a98: color = 2'b11;
      13'h1a99: color = 2'b11;
      13'h1a9a: color = 2'b00;
      13'h1a9b: color = 2'b00;
      13'h1a9c: color = 2'b10;
      13'h1a9d: color = 2'b10;
      13'h1a9e: color = 2'b11;
      13'h1a9f: color = 2'b11;
      13'h1aa0: color = 2'b10;
      13'h1aa1: color = 2'b10;
      13'h1aa2: color = 2'b00;
      13'h1aa3: color = 2'b00;
      13'h1aa4: color = 2'b00;
      13'h1aa5: color = 2'b00;
      13'h1aa6: color = 2'b00;
      13'h1aa7: color = 2'b00;
      13'h1aa8: color = 2'b00;
      13'h1aa9: color = 2'b00;
      13'h1aaa: color = 2'b00;
      13'h1aab: color = 2'b00;
      13'h1aac: color = 2'b00;
      13'h1aad: color = 2'b00;
      13'h1aae: color = 2'b00;
      13'h1aaf: color = 2'b00;
      13'h1ab0: color = 2'b00;
      13'h1ab1: color = 2'b00;
      13'h1ab2: color = 2'b00;
      13'h1ab3: color = 2'b00;
      13'h1ab4: color = 2'b00;
      13'h1ab5: color = 2'b00;
      13'h1ab6: color = 2'b00;
      13'h1ab7: color = 2'b00;
      13'h1ab8: color = 2'b00;
      13'h1ab9: color = 2'b00;
      13'h1aba: color = 2'b00;
      13'h1abb: color = 2'b00;
      13'h1abc: color = 2'b00;
      13'h1abd: color = 2'b00;
      13'h1abe: color = 2'b00;
      13'h1abf: color = 2'b00;
      13'h1ac0: color = 2'b00;
      13'h1ac1: color = 2'b00;
      13'h1ac2: color = 2'b00;
      13'h1ac3: color = 2'b00;
      13'h1ac4: color = 2'b00;
      13'h1ac5: color = 2'b00;
      13'h1ac6: color = 2'b00;
      13'h1ac7: color = 2'b00;
      13'h1ac8: color = 2'b00;
      13'h1ac9: color = 2'b00;
      13'h1aca: color = 2'b00;
      13'h1acb: color = 2'b00;
      13'h1acc: color = 2'b00;
      13'h1acd: color = 2'b00;
      13'h1ace: color = 2'b00;
      13'h1acf: color = 2'b00;
      13'h1ad0: color = 2'b00;
      13'h1ad1: color = 2'b00;
      13'h1ad2: color = 2'b00;
      13'h1ad3: color = 2'b00;
      13'h1ad4: color = 2'b00;
      13'h1ad5: color = 2'b00;
      13'h1ad6: color = 2'b00;
      13'h1ad7: color = 2'b00;
      13'h1ad8: color = 2'b00;
      13'h1ad9: color = 2'b00;
      13'h1ada: color = 2'b00;
      13'h1adb: color = 2'b00;
      13'h1adc: color = 2'b00;
      13'h1add: color = 2'b00;
      13'h1ade: color = 2'b11;
      13'h1adf: color = 2'b11;
      13'h1ae0: color = 2'b10;
      13'h1ae1: color = 2'b10;
      13'h1ae2: color = 2'b11;
      13'h1ae3: color = 2'b11;
      13'h1ae4: color = 2'b00;
      13'h1ae5: color = 2'b00;
      13'h1ae6: color = 2'b11;
      13'h1ae7: color = 2'b11;
      13'h1ae8: color = 2'b11;
      13'h1ae9: color = 2'b11;
      13'h1aea: color = 2'b11;
      13'h1aeb: color = 2'b11;
      13'h1aec: color = 2'b11;
      13'h1aed: color = 2'b11;
      13'h1aee: color = 2'b11;
      13'h1aef: color = 2'b11;
      13'h1af0: color = 2'b11;
      13'h1af1: color = 2'b11;
      13'h1af2: color = 2'b11;
      13'h1af3: color = 2'b11;
      13'h1af4: color = 2'b11;
      13'h1af5: color = 2'b11;
      13'h1af6: color = 2'b11;
      13'h1af7: color = 2'b11;
      13'h1af8: color = 2'b11;
      13'h1af9: color = 2'b11;
      13'h1afa: color = 2'b00;
      13'h1afb: color = 2'b00;
      13'h1afc: color = 2'b10;
      13'h1afd: color = 2'b10;
      13'h1afe: color = 2'b11;
      13'h1aff: color = 2'b11;
      13'h1b00: color = 2'b11;
      13'h1b01: color = 2'b11;
      13'h1b02: color = 2'b11;
      13'h1b03: color = 2'b11;
      13'h1b04: color = 2'b00;
      13'h1b05: color = 2'b00;
      13'h1b06: color = 2'b10;
      13'h1b07: color = 2'b10;
      13'h1b08: color = 2'b10;
      13'h1b09: color = 2'b10;
      13'h1b0a: color = 2'b10;
      13'h1b0b: color = 2'b10;
      13'h1b0c: color = 2'b10;
      13'h1b0d: color = 2'b10;
      13'h1b0e: color = 2'b10;
      13'h1b0f: color = 2'b10;
      13'h1b10: color = 2'b10;
      13'h1b11: color = 2'b10;
      13'h1b12: color = 2'b10;
      13'h1b13: color = 2'b10;
      13'h1b14: color = 2'b10;
      13'h1b15: color = 2'b10;
      13'h1b16: color = 2'b10;
      13'h1b17: color = 2'b10;
      13'h1b18: color = 2'b10;
      13'h1b19: color = 2'b10;
      13'h1b1a: color = 2'b00;
      13'h1b1b: color = 2'b00;
      13'h1b1c: color = 2'b11;
      13'h1b1d: color = 2'b11;
      13'h1b1e: color = 2'b10;
      13'h1b1f: color = 2'b10;
      13'h1b20: color = 2'b11;
      13'h1b21: color = 2'b11;
      13'h1b22: color = 2'b00;
      13'h1b23: color = 2'b00;
      13'h1b24: color = 2'b01;
      13'h1b25: color = 2'b01;
      13'h1b26: color = 2'b01;
      13'h1b27: color = 2'b01;
      13'h1b28: color = 2'b01;
      13'h1b29: color = 2'b01;
      13'h1b2a: color = 2'b00;
      13'h1b2b: color = 2'b00;
      13'h1b2c: color = 2'b01;
      13'h1b2d: color = 2'b01;
      13'h1b2e: color = 2'b01;
      13'h1b2f: color = 2'b01;
      13'h1b30: color = 2'b01;
      13'h1b31: color = 2'b01;
      13'h1b32: color = 2'b01;
      13'h1b33: color = 2'b01;
      13'h1b34: color = 2'b01;
      13'h1b35: color = 2'b01;
      13'h1b36: color = 2'b01;
      13'h1b37: color = 2'b01;
      13'h1b38: color = 2'b01;
      13'h1b39: color = 2'b01;
      13'h1b3a: color = 2'b01;
      13'h1b3b: color = 2'b01;
      13'h1b3c: color = 2'b01;
      13'h1b3d: color = 2'b01;
      13'h1b3e: color = 2'b01;
      13'h1b3f: color = 2'b01;
      13'h1b40: color = 2'b01;
      13'h1b41: color = 2'b01;
      13'h1b42: color = 2'b01;
      13'h1b43: color = 2'b01;
      13'h1b44: color = 2'b01;
      13'h1b45: color = 2'b01;
      13'h1b46: color = 2'b01;
      13'h1b47: color = 2'b01;
      13'h1b48: color = 2'b01;
      13'h1b49: color = 2'b01;
      13'h1b4a: color = 2'b01;
      13'h1b4b: color = 2'b01;
      13'h1b4c: color = 2'b01;
      13'h1b4d: color = 2'b01;
      13'h1b4e: color = 2'b01;
      13'h1b4f: color = 2'b01;
      13'h1b50: color = 2'b01;
      13'h1b51: color = 2'b01;
      13'h1b52: color = 2'b01;
      13'h1b53: color = 2'b01;
      13'h1b54: color = 2'b00;
      13'h1b55: color = 2'b00;
      13'h1b56: color = 2'b01;
      13'h1b57: color = 2'b01;
      13'h1b58: color = 2'b01;
      13'h1b59: color = 2'b01;
      13'h1b5a: color = 2'b01;
      13'h1b5b: color = 2'b01;
      13'h1b5c: color = 2'b00;
      13'h1b5d: color = 2'b00;
      13'h1b5e: color = 2'b10;
      13'h1b5f: color = 2'b10;
      13'h1b60: color = 2'b11;
      13'h1b61: color = 2'b11;
      13'h1b62: color = 2'b11;
      13'h1b63: color = 2'b11;
      13'h1b64: color = 2'b00;
      13'h1b65: color = 2'b00;
      13'h1b66: color = 2'b10;
      13'h1b67: color = 2'b10;
      13'h1b68: color = 2'b10;
      13'h1b69: color = 2'b10;
      13'h1b6a: color = 2'b10;
      13'h1b6b: color = 2'b10;
      13'h1b6c: color = 2'b10;
      13'h1b6d: color = 2'b10;
      13'h1b6e: color = 2'b10;
      13'h1b6f: color = 2'b10;
      13'h1b70: color = 2'b10;
      13'h1b71: color = 2'b10;
      13'h1b72: color = 2'b10;
      13'h1b73: color = 2'b10;
      13'h1b74: color = 2'b10;
      13'h1b75: color = 2'b10;
      13'h1b76: color = 2'b10;
      13'h1b77: color = 2'b10;
      13'h1b78: color = 2'b10;
      13'h1b79: color = 2'b10;
      13'h1b7a: color = 2'b00;
      13'h1b7b: color = 2'b00;
      13'h1b7c: color = 2'b11;
      13'h1b7d: color = 2'b11;
      13'h1b7e: color = 2'b10;
      13'h1b7f: color = 2'b10;
      13'h1b80: color = 2'b11;
      13'h1b81: color = 2'b11;
      13'h1b82: color = 2'b11;
      13'h1b83: color = 2'b11;
      13'h1b84: color = 2'b00;
      13'h1b85: color = 2'b00;
      13'h1b86: color = 2'b10;
      13'h1b87: color = 2'b10;
      13'h1b88: color = 2'b10;
      13'h1b89: color = 2'b10;
      13'h1b8a: color = 2'b10;
      13'h1b8b: color = 2'b10;
      13'h1b8c: color = 2'b10;
      13'h1b8d: color = 2'b10;
      13'h1b8e: color = 2'b10;
      13'h1b8f: color = 2'b10;
      13'h1b90: color = 2'b10;
      13'h1b91: color = 2'b10;
      13'h1b92: color = 2'b10;
      13'h1b93: color = 2'b10;
      13'h1b94: color = 2'b10;
      13'h1b95: color = 2'b10;
      13'h1b96: color = 2'b10;
      13'h1b97: color = 2'b10;
      13'h1b98: color = 2'b10;
      13'h1b99: color = 2'b10;
      13'h1b9a: color = 2'b00;
      13'h1b9b: color = 2'b00;
      13'h1b9c: color = 2'b11;
      13'h1b9d: color = 2'b11;
      13'h1b9e: color = 2'b10;
      13'h1b9f: color = 2'b10;
      13'h1ba0: color = 2'b11;
      13'h1ba1: color = 2'b11;
      13'h1ba2: color = 2'b00;
      13'h1ba3: color = 2'b00;
      13'h1ba4: color = 2'b01;
      13'h1ba5: color = 2'b01;
      13'h1ba6: color = 2'b01;
      13'h1ba7: color = 2'b01;
      13'h1ba8: color = 2'b01;
      13'h1ba9: color = 2'b01;
      13'h1baa: color = 2'b00;
      13'h1bab: color = 2'b00;
      13'h1bac: color = 2'b01;
      13'h1bad: color = 2'b01;
      13'h1bae: color = 2'b01;
      13'h1baf: color = 2'b01;
      13'h1bb0: color = 2'b01;
      13'h1bb1: color = 2'b01;
      13'h1bb2: color = 2'b01;
      13'h1bb3: color = 2'b01;
      13'h1bb4: color = 2'b01;
      13'h1bb5: color = 2'b01;
      13'h1bb6: color = 2'b01;
      13'h1bb7: color = 2'b01;
      13'h1bb8: color = 2'b01;
      13'h1bb9: color = 2'b01;
      13'h1bba: color = 2'b01;
      13'h1bbb: color = 2'b01;
      13'h1bbc: color = 2'b01;
      13'h1bbd: color = 2'b01;
      13'h1bbe: color = 2'b01;
      13'h1bbf: color = 2'b01;
      13'h1bc0: color = 2'b01;
      13'h1bc1: color = 2'b01;
      13'h1bc2: color = 2'b01;
      13'h1bc3: color = 2'b01;
      13'h1bc4: color = 2'b01;
      13'h1bc5: color = 2'b01;
      13'h1bc6: color = 2'b01;
      13'h1bc7: color = 2'b01;
      13'h1bc8: color = 2'b01;
      13'h1bc9: color = 2'b01;
      13'h1bca: color = 2'b01;
      13'h1bcb: color = 2'b01;
      13'h1bcc: color = 2'b01;
      13'h1bcd: color = 2'b01;
      13'h1bce: color = 2'b01;
      13'h1bcf: color = 2'b01;
      13'h1bd0: color = 2'b01;
      13'h1bd1: color = 2'b01;
      13'h1bd2: color = 2'b01;
      13'h1bd3: color = 2'b01;
      13'h1bd4: color = 2'b00;
      13'h1bd5: color = 2'b00;
      13'h1bd6: color = 2'b01;
      13'h1bd7: color = 2'b01;
      13'h1bd8: color = 2'b01;
      13'h1bd9: color = 2'b01;
      13'h1bda: color = 2'b01;
      13'h1bdb: color = 2'b01;
      13'h1bdc: color = 2'b00;
      13'h1bdd: color = 2'b00;
      13'h1bde: color = 2'b10;
      13'h1bdf: color = 2'b10;
      13'h1be0: color = 2'b11;
      13'h1be1: color = 2'b11;
      13'h1be2: color = 2'b11;
      13'h1be3: color = 2'b11;
      13'h1be4: color = 2'b00;
      13'h1be5: color = 2'b00;
      13'h1be6: color = 2'b10;
      13'h1be7: color = 2'b10;
      13'h1be8: color = 2'b10;
      13'h1be9: color = 2'b10;
      13'h1bea: color = 2'b10;
      13'h1beb: color = 2'b10;
      13'h1bec: color = 2'b10;
      13'h1bed: color = 2'b10;
      13'h1bee: color = 2'b10;
      13'h1bef: color = 2'b10;
      13'h1bf0: color = 2'b10;
      13'h1bf1: color = 2'b10;
      13'h1bf2: color = 2'b10;
      13'h1bf3: color = 2'b10;
      13'h1bf4: color = 2'b10;
      13'h1bf5: color = 2'b10;
      13'h1bf6: color = 2'b10;
      13'h1bf7: color = 2'b10;
      13'h1bf8: color = 2'b10;
      13'h1bf9: color = 2'b10;
      13'h1bfa: color = 2'b00;
      13'h1bfb: color = 2'b00;
      13'h1bfc: color = 2'b11;
      13'h1bfd: color = 2'b11;
      13'h1bfe: color = 2'b10;
      13'h1bff: color = 2'b10;
      13'h1c00: color = 2'b10;
      13'h1c01: color = 2'b10;
      13'h1c02: color = 2'b11;
      13'h1c03: color = 2'b11;
      13'h1c04: color = 2'b00;
      13'h1c05: color = 2'b00;
      13'h1c06: color = 2'b10;
      13'h1c07: color = 2'b10;
      13'h1c08: color = 2'b00;
      13'h1c09: color = 2'b00;
      13'h1c0a: color = 2'b00;
      13'h1c0b: color = 2'b00;
      13'h1c0c: color = 2'b00;
      13'h1c0d: color = 2'b00;
      13'h1c0e: color = 2'b00;
      13'h1c0f: color = 2'b00;
      13'h1c10: color = 2'b00;
      13'h1c11: color = 2'b00;
      13'h1c12: color = 2'b00;
      13'h1c13: color = 2'b00;
      13'h1c14: color = 2'b00;
      13'h1c15: color = 2'b00;
      13'h1c16: color = 2'b00;
      13'h1c17: color = 2'b00;
      13'h1c18: color = 2'b10;
      13'h1c19: color = 2'b10;
      13'h1c1a: color = 2'b00;
      13'h1c1b: color = 2'b00;
      13'h1c1c: color = 2'b11;
      13'h1c1d: color = 2'b11;
      13'h1c1e: color = 2'b11;
      13'h1c1f: color = 2'b11;
      13'h1c20: color = 2'b10;
      13'h1c21: color = 2'b10;
      13'h1c22: color = 2'b00;
      13'h1c23: color = 2'b00;
      13'h1c24: color = 2'b11;
      13'h1c25: color = 2'b11;
      13'h1c26: color = 2'b10;
      13'h1c27: color = 2'b10;
      13'h1c28: color = 2'b10;
      13'h1c29: color = 2'b10;
      13'h1c2a: color = 2'b00;
      13'h1c2b: color = 2'b00;
      13'h1c2c: color = 2'b00;
      13'h1c2d: color = 2'b00;
      13'h1c2e: color = 2'b00;
      13'h1c2f: color = 2'b00;
      13'h1c30: color = 2'b00;
      13'h1c31: color = 2'b00;
      13'h1c32: color = 2'b00;
      13'h1c33: color = 2'b00;
      13'h1c34: color = 2'b00;
      13'h1c35: color = 2'b00;
      13'h1c36: color = 2'b00;
      13'h1c37: color = 2'b00;
      13'h1c38: color = 2'b00;
      13'h1c39: color = 2'b00;
      13'h1c3a: color = 2'b00;
      13'h1c3b: color = 2'b00;
      13'h1c3c: color = 2'b00;
      13'h1c3d: color = 2'b00;
      13'h1c3e: color = 2'b00;
      13'h1c3f: color = 2'b00;
      13'h1c40: color = 2'b00;
      13'h1c41: color = 2'b00;
      13'h1c42: color = 2'b00;
      13'h1c43: color = 2'b00;
      13'h1c44: color = 2'b00;
      13'h1c45: color = 2'b00;
      13'h1c46: color = 2'b00;
      13'h1c47: color = 2'b00;
      13'h1c48: color = 2'b00;
      13'h1c49: color = 2'b00;
      13'h1c4a: color = 2'b00;
      13'h1c4b: color = 2'b00;
      13'h1c4c: color = 2'b00;
      13'h1c4d: color = 2'b00;
      13'h1c4e: color = 2'b00;
      13'h1c4f: color = 2'b00;
      13'h1c50: color = 2'b00;
      13'h1c51: color = 2'b00;
      13'h1c52: color = 2'b00;
      13'h1c53: color = 2'b00;
      13'h1c54: color = 2'b00;
      13'h1c55: color = 2'b00;
      13'h1c56: color = 2'b10;
      13'h1c57: color = 2'b10;
      13'h1c58: color = 2'b10;
      13'h1c59: color = 2'b10;
      13'h1c5a: color = 2'b10;
      13'h1c5b: color = 2'b10;
      13'h1c5c: color = 2'b00;
      13'h1c5d: color = 2'b00;
      13'h1c5e: color = 2'b11;
      13'h1c5f: color = 2'b11;
      13'h1c60: color = 2'b10;
      13'h1c61: color = 2'b10;
      13'h1c62: color = 2'b11;
      13'h1c63: color = 2'b11;
      13'h1c64: color = 2'b00;
      13'h1c65: color = 2'b00;
      13'h1c66: color = 2'b10;
      13'h1c67: color = 2'b10;
      13'h1c68: color = 2'b00;
      13'h1c69: color = 2'b00;
      13'h1c6a: color = 2'b00;
      13'h1c6b: color = 2'b00;
      13'h1c6c: color = 2'b00;
      13'h1c6d: color = 2'b00;
      13'h1c6e: color = 2'b00;
      13'h1c6f: color = 2'b00;
      13'h1c70: color = 2'b00;
      13'h1c71: color = 2'b00;
      13'h1c72: color = 2'b00;
      13'h1c73: color = 2'b00;
      13'h1c74: color = 2'b00;
      13'h1c75: color = 2'b00;
      13'h1c76: color = 2'b00;
      13'h1c77: color = 2'b00;
      13'h1c78: color = 2'b10;
      13'h1c79: color = 2'b10;
      13'h1c7a: color = 2'b00;
      13'h1c7b: color = 2'b00;
      13'h1c7c: color = 2'b11;
      13'h1c7d: color = 2'b11;
      13'h1c7e: color = 2'b11;
      13'h1c7f: color = 2'b11;
      13'h1c80: color = 2'b10;
      13'h1c81: color = 2'b10;
      13'h1c82: color = 2'b11;
      13'h1c83: color = 2'b11;
      13'h1c84: color = 2'b00;
      13'h1c85: color = 2'b00;
      13'h1c86: color = 2'b10;
      13'h1c87: color = 2'b10;
      13'h1c88: color = 2'b00;
      13'h1c89: color = 2'b00;
      13'h1c8a: color = 2'b00;
      13'h1c8b: color = 2'b00;
      13'h1c8c: color = 2'b00;
      13'h1c8d: color = 2'b00;
      13'h1c8e: color = 2'b00;
      13'h1c8f: color = 2'b00;
      13'h1c90: color = 2'b00;
      13'h1c91: color = 2'b00;
      13'h1c92: color = 2'b00;
      13'h1c93: color = 2'b00;
      13'h1c94: color = 2'b00;
      13'h1c95: color = 2'b00;
      13'h1c96: color = 2'b00;
      13'h1c97: color = 2'b00;
      13'h1c98: color = 2'b10;
      13'h1c99: color = 2'b10;
      13'h1c9a: color = 2'b00;
      13'h1c9b: color = 2'b00;
      13'h1c9c: color = 2'b11;
      13'h1c9d: color = 2'b11;
      13'h1c9e: color = 2'b11;
      13'h1c9f: color = 2'b11;
      13'h1ca0: color = 2'b10;
      13'h1ca1: color = 2'b10;
      13'h1ca2: color = 2'b00;
      13'h1ca3: color = 2'b00;
      13'h1ca4: color = 2'b11;
      13'h1ca5: color = 2'b11;
      13'h1ca6: color = 2'b10;
      13'h1ca7: color = 2'b10;
      13'h1ca8: color = 2'b10;
      13'h1ca9: color = 2'b10;
      13'h1caa: color = 2'b00;
      13'h1cab: color = 2'b00;
      13'h1cac: color = 2'b00;
      13'h1cad: color = 2'b00;
      13'h1cae: color = 2'b00;
      13'h1caf: color = 2'b00;
      13'h1cb0: color = 2'b00;
      13'h1cb1: color = 2'b00;
      13'h1cb2: color = 2'b00;
      13'h1cb3: color = 2'b00;
      13'h1cb4: color = 2'b00;
      13'h1cb5: color = 2'b00;
      13'h1cb6: color = 2'b00;
      13'h1cb7: color = 2'b00;
      13'h1cb8: color = 2'b00;
      13'h1cb9: color = 2'b00;
      13'h1cba: color = 2'b00;
      13'h1cbb: color = 2'b00;
      13'h1cbc: color = 2'b00;
      13'h1cbd: color = 2'b00;
      13'h1cbe: color = 2'b00;
      13'h1cbf: color = 2'b00;
      13'h1cc0: color = 2'b00;
      13'h1cc1: color = 2'b00;
      13'h1cc2: color = 2'b00;
      13'h1cc3: color = 2'b00;
      13'h1cc4: color = 2'b00;
      13'h1cc5: color = 2'b00;
      13'h1cc6: color = 2'b00;
      13'h1cc7: color = 2'b00;
      13'h1cc8: color = 2'b00;
      13'h1cc9: color = 2'b00;
      13'h1cca: color = 2'b00;
      13'h1ccb: color = 2'b00;
      13'h1ccc: color = 2'b00;
      13'h1ccd: color = 2'b00;
      13'h1cce: color = 2'b00;
      13'h1ccf: color = 2'b00;
      13'h1cd0: color = 2'b00;
      13'h1cd1: color = 2'b00;
      13'h1cd2: color = 2'b00;
      13'h1cd3: color = 2'b00;
      13'h1cd4: color = 2'b00;
      13'h1cd5: color = 2'b00;
      13'h1cd6: color = 2'b10;
      13'h1cd7: color = 2'b10;
      13'h1cd8: color = 2'b10;
      13'h1cd9: color = 2'b10;
      13'h1cda: color = 2'b10;
      13'h1cdb: color = 2'b10;
      13'h1cdc: color = 2'b00;
      13'h1cdd: color = 2'b00;
      13'h1cde: color = 2'b11;
      13'h1cdf: color = 2'b11;
      13'h1ce0: color = 2'b10;
      13'h1ce1: color = 2'b10;
      13'h1ce2: color = 2'b11;
      13'h1ce3: color = 2'b11;
      13'h1ce4: color = 2'b00;
      13'h1ce5: color = 2'b00;
      13'h1ce6: color = 2'b10;
      13'h1ce7: color = 2'b10;
      13'h1ce8: color = 2'b00;
      13'h1ce9: color = 2'b00;
      13'h1cea: color = 2'b00;
      13'h1ceb: color = 2'b00;
      13'h1cec: color = 2'b00;
      13'h1ced: color = 2'b00;
      13'h1cee: color = 2'b00;
      13'h1cef: color = 2'b00;
      13'h1cf0: color = 2'b00;
      13'h1cf1: color = 2'b00;
      13'h1cf2: color = 2'b00;
      13'h1cf3: color = 2'b00;
      13'h1cf4: color = 2'b00;
      13'h1cf5: color = 2'b00;
      13'h1cf6: color = 2'b00;
      13'h1cf7: color = 2'b00;
      13'h1cf8: color = 2'b10;
      13'h1cf9: color = 2'b10;
      13'h1cfa: color = 2'b00;
      13'h1cfb: color = 2'b00;
      13'h1cfc: color = 2'b11;
      13'h1cfd: color = 2'b11;
      13'h1cfe: color = 2'b11;
      13'h1cff: color = 2'b11;
      13'h1d00: color = 2'b11;
      13'h1d01: color = 2'b11;
      13'h1d02: color = 2'b10;
      13'h1d03: color = 2'b10;
      13'h1d04: color = 2'b00;
      13'h1d05: color = 2'b00;
      13'h1d06: color = 2'b10;
      13'h1d07: color = 2'b10;
      13'h1d08: color = 2'b00;
      13'h1d09: color = 2'b00;
      13'h1d0a: color = 2'b11;
      13'h1d0b: color = 2'b11;
      13'h1d0c: color = 2'b11;
      13'h1d0d: color = 2'b11;
      13'h1d0e: color = 2'b11;
      13'h1d0f: color = 2'b11;
      13'h1d10: color = 2'b11;
      13'h1d11: color = 2'b11;
      13'h1d12: color = 2'b10;
      13'h1d13: color = 2'b10;
      13'h1d14: color = 2'b11;
      13'h1d15: color = 2'b11;
      13'h1d16: color = 2'b00;
      13'h1d17: color = 2'b00;
      13'h1d18: color = 2'b10;
      13'h1d19: color = 2'b10;
      13'h1d1a: color = 2'b00;
      13'h1d1b: color = 2'b00;
      13'h1d1c: color = 2'b11;
      13'h1d1d: color = 2'b11;
      13'h1d1e: color = 2'b11;
      13'h1d1f: color = 2'b11;
      13'h1d20: color = 2'b11;
      13'h1d21: color = 2'b11;
      13'h1d22: color = 2'b00;
      13'h1d23: color = 2'b00;
      13'h1d24: color = 2'b11;
      13'h1d25: color = 2'b11;
      13'h1d26: color = 2'b10;
      13'h1d27: color = 2'b10;
      13'h1d28: color = 2'b10;
      13'h1d29: color = 2'b10;
      13'h1d2a: color = 2'b00;
      13'h1d2b: color = 2'b00;
      13'h1d2c: color = 2'b10;
      13'h1d2d: color = 2'b10;
      13'h1d2e: color = 2'b10;
      13'h1d2f: color = 2'b10;
      13'h1d30: color = 2'b10;
      13'h1d31: color = 2'b10;
      13'h1d32: color = 2'b10;
      13'h1d33: color = 2'b10;
      13'h1d34: color = 2'b10;
      13'h1d35: color = 2'b10;
      13'h1d36: color = 2'b10;
      13'h1d37: color = 2'b10;
      13'h1d38: color = 2'b10;
      13'h1d39: color = 2'b10;
      13'h1d3a: color = 2'b10;
      13'h1d3b: color = 2'b10;
      13'h1d3c: color = 2'b10;
      13'h1d3d: color = 2'b10;
      13'h1d3e: color = 2'b10;
      13'h1d3f: color = 2'b10;
      13'h1d40: color = 2'b10;
      13'h1d41: color = 2'b10;
      13'h1d42: color = 2'b10;
      13'h1d43: color = 2'b10;
      13'h1d44: color = 2'b10;
      13'h1d45: color = 2'b10;
      13'h1d46: color = 2'b10;
      13'h1d47: color = 2'b10;
      13'h1d48: color = 2'b10;
      13'h1d49: color = 2'b10;
      13'h1d4a: color = 2'b10;
      13'h1d4b: color = 2'b10;
      13'h1d4c: color = 2'b10;
      13'h1d4d: color = 2'b10;
      13'h1d4e: color = 2'b10;
      13'h1d4f: color = 2'b10;
      13'h1d50: color = 2'b10;
      13'h1d51: color = 2'b10;
      13'h1d52: color = 2'b10;
      13'h1d53: color = 2'b10;
      13'h1d54: color = 2'b00;
      13'h1d55: color = 2'b00;
      13'h1d56: color = 2'b10;
      13'h1d57: color = 2'b10;
      13'h1d58: color = 2'b10;
      13'h1d59: color = 2'b10;
      13'h1d5a: color = 2'b10;
      13'h1d5b: color = 2'b10;
      13'h1d5c: color = 2'b00;
      13'h1d5d: color = 2'b00;
      13'h1d5e: color = 2'b11;
      13'h1d5f: color = 2'b11;
      13'h1d60: color = 2'b11;
      13'h1d61: color = 2'b11;
      13'h1d62: color = 2'b10;
      13'h1d63: color = 2'b10;
      13'h1d64: color = 2'b00;
      13'h1d65: color = 2'b00;
      13'h1d66: color = 2'b10;
      13'h1d67: color = 2'b10;
      13'h1d68: color = 2'b00;
      13'h1d69: color = 2'b00;
      13'h1d6a: color = 2'b11;
      13'h1d6b: color = 2'b11;
      13'h1d6c: color = 2'b11;
      13'h1d6d: color = 2'b11;
      13'h1d6e: color = 2'b11;
      13'h1d6f: color = 2'b11;
      13'h1d70: color = 2'b11;
      13'h1d71: color = 2'b11;
      13'h1d72: color = 2'b10;
      13'h1d73: color = 2'b10;
      13'h1d74: color = 2'b11;
      13'h1d75: color = 2'b11;
      13'h1d76: color = 2'b00;
      13'h1d77: color = 2'b00;
      13'h1d78: color = 2'b10;
      13'h1d79: color = 2'b10;
      13'h1d7a: color = 2'b00;
      13'h1d7b: color = 2'b00;
      13'h1d7c: color = 2'b11;
      13'h1d7d: color = 2'b11;
      13'h1d7e: color = 2'b11;
      13'h1d7f: color = 2'b11;
      13'h1d80: color = 2'b11;
      13'h1d81: color = 2'b11;
      13'h1d82: color = 2'b10;
      13'h1d83: color = 2'b10;
      13'h1d84: color = 2'b00;
      13'h1d85: color = 2'b00;
      13'h1d86: color = 2'b10;
      13'h1d87: color = 2'b10;
      13'h1d88: color = 2'b00;
      13'h1d89: color = 2'b00;
      13'h1d8a: color = 2'b11;
      13'h1d8b: color = 2'b11;
      13'h1d8c: color = 2'b11;
      13'h1d8d: color = 2'b11;
      13'h1d8e: color = 2'b11;
      13'h1d8f: color = 2'b11;
      13'h1d90: color = 2'b11;
      13'h1d91: color = 2'b11;
      13'h1d92: color = 2'b10;
      13'h1d93: color = 2'b10;
      13'h1d94: color = 2'b11;
      13'h1d95: color = 2'b11;
      13'h1d96: color = 2'b00;
      13'h1d97: color = 2'b00;
      13'h1d98: color = 2'b10;
      13'h1d99: color = 2'b10;
      13'h1d9a: color = 2'b00;
      13'h1d9b: color = 2'b00;
      13'h1d9c: color = 2'b11;
      13'h1d9d: color = 2'b11;
      13'h1d9e: color = 2'b11;
      13'h1d9f: color = 2'b11;
      13'h1da0: color = 2'b11;
      13'h1da1: color = 2'b11;
      13'h1da2: color = 2'b00;
      13'h1da3: color = 2'b00;
      13'h1da4: color = 2'b11;
      13'h1da5: color = 2'b11;
      13'h1da6: color = 2'b10;
      13'h1da7: color = 2'b10;
      13'h1da8: color = 2'b10;
      13'h1da9: color = 2'b10;
      13'h1daa: color = 2'b00;
      13'h1dab: color = 2'b00;
      13'h1dac: color = 2'b10;
      13'h1dad: color = 2'b10;
      13'h1dae: color = 2'b10;
      13'h1daf: color = 2'b10;
      13'h1db0: color = 2'b10;
      13'h1db1: color = 2'b10;
      13'h1db2: color = 2'b10;
      13'h1db3: color = 2'b10;
      13'h1db4: color = 2'b10;
      13'h1db5: color = 2'b10;
      13'h1db6: color = 2'b10;
      13'h1db7: color = 2'b10;
      13'h1db8: color = 2'b10;
      13'h1db9: color = 2'b10;
      13'h1dba: color = 2'b10;
      13'h1dbb: color = 2'b10;
      13'h1dbc: color = 2'b10;
      13'h1dbd: color = 2'b10;
      13'h1dbe: color = 2'b10;
      13'h1dbf: color = 2'b10;
      13'h1dc0: color = 2'b10;
      13'h1dc1: color = 2'b10;
      13'h1dc2: color = 2'b10;
      13'h1dc3: color = 2'b10;
      13'h1dc4: color = 2'b10;
      13'h1dc5: color = 2'b10;
      13'h1dc6: color = 2'b10;
      13'h1dc7: color = 2'b10;
      13'h1dc8: color = 2'b10;
      13'h1dc9: color = 2'b10;
      13'h1dca: color = 2'b10;
      13'h1dcb: color = 2'b10;
      13'h1dcc: color = 2'b10;
      13'h1dcd: color = 2'b10;
      13'h1dce: color = 2'b10;
      13'h1dcf: color = 2'b10;
      13'h1dd0: color = 2'b10;
      13'h1dd1: color = 2'b10;
      13'h1dd2: color = 2'b10;
      13'h1dd3: color = 2'b10;
      13'h1dd4: color = 2'b00;
      13'h1dd5: color = 2'b00;
      13'h1dd6: color = 2'b10;
      13'h1dd7: color = 2'b10;
      13'h1dd8: color = 2'b10;
      13'h1dd9: color = 2'b10;
      13'h1dda: color = 2'b10;
      13'h1ddb: color = 2'b10;
      13'h1ddc: color = 2'b00;
      13'h1ddd: color = 2'b00;
      13'h1dde: color = 2'b11;
      13'h1ddf: color = 2'b11;
      13'h1de0: color = 2'b11;
      13'h1de1: color = 2'b11;
      13'h1de2: color = 2'b10;
      13'h1de3: color = 2'b10;
      13'h1de4: color = 2'b00;
      13'h1de5: color = 2'b00;
      13'h1de6: color = 2'b10;
      13'h1de7: color = 2'b10;
      13'h1de8: color = 2'b00;
      13'h1de9: color = 2'b00;
      13'h1dea: color = 2'b11;
      13'h1deb: color = 2'b11;
      13'h1dec: color = 2'b11;
      13'h1ded: color = 2'b11;
      13'h1dee: color = 2'b11;
      13'h1def: color = 2'b11;
      13'h1df0: color = 2'b11;
      13'h1df1: color = 2'b11;
      13'h1df2: color = 2'b10;
      13'h1df3: color = 2'b10;
      13'h1df4: color = 2'b11;
      13'h1df5: color = 2'b11;
      13'h1df6: color = 2'b00;
      13'h1df7: color = 2'b00;
      13'h1df8: color = 2'b10;
      13'h1df9: color = 2'b10;
      13'h1dfa: color = 2'b00;
      13'h1dfb: color = 2'b00;
      13'h1dfc: color = 2'b11;
      13'h1dfd: color = 2'b11;
      13'h1dfe: color = 2'b11;
      13'h1dff: color = 2'b11;
      13'h1e00: color = 2'b11;
      13'h1e01: color = 2'b11;
      13'h1e02: color = 2'b11;
      13'h1e03: color = 2'b11;
      13'h1e04: color = 2'b00;
      13'h1e05: color = 2'b00;
      13'h1e06: color = 2'b10;
      13'h1e07: color = 2'b10;
      13'h1e08: color = 2'b00;
      13'h1e09: color = 2'b00;
      13'h1e0a: color = 2'b11;
      13'h1e0b: color = 2'b11;
      13'h1e0c: color = 2'b11;
      13'h1e0d: color = 2'b11;
      13'h1e0e: color = 2'b11;
      13'h1e0f: color = 2'b11;
      13'h1e10: color = 2'b11;
      13'h1e11: color = 2'b11;
      13'h1e12: color = 2'b11;
      13'h1e13: color = 2'b11;
      13'h1e14: color = 2'b10;
      13'h1e15: color = 2'b10;
      13'h1e16: color = 2'b00;
      13'h1e17: color = 2'b00;
      13'h1e18: color = 2'b10;
      13'h1e19: color = 2'b10;
      13'h1e1a: color = 2'b00;
      13'h1e1b: color = 2'b00;
      13'h1e1c: color = 2'b11;
      13'h1e1d: color = 2'b11;
      13'h1e1e: color = 2'b11;
      13'h1e1f: color = 2'b11;
      13'h1e20: color = 2'b11;
      13'h1e21: color = 2'b11;
      13'h1e22: color = 2'b00;
      13'h1e23: color = 2'b00;
      13'h1e24: color = 2'b00;
      13'h1e25: color = 2'b00;
      13'h1e26: color = 2'b00;
      13'h1e27: color = 2'b00;
      13'h1e28: color = 2'b00;
      13'h1e29: color = 2'b00;
      13'h1e2a: color = 2'b00;
      13'h1e2b: color = 2'b00;
      13'h1e2c: color = 2'b10;
      13'h1e2d: color = 2'b10;
      13'h1e2e: color = 2'b10;
      13'h1e2f: color = 2'b10;
      13'h1e30: color = 2'b10;
      13'h1e31: color = 2'b10;
      13'h1e32: color = 2'b10;
      13'h1e33: color = 2'b10;
      13'h1e34: color = 2'b10;
      13'h1e35: color = 2'b10;
      13'h1e36: color = 2'b10;
      13'h1e37: color = 2'b10;
      13'h1e38: color = 2'b10;
      13'h1e39: color = 2'b10;
      13'h1e3a: color = 2'b10;
      13'h1e3b: color = 2'b10;
      13'h1e3c: color = 2'b10;
      13'h1e3d: color = 2'b10;
      13'h1e3e: color = 2'b10;
      13'h1e3f: color = 2'b10;
      13'h1e40: color = 2'b10;
      13'h1e41: color = 2'b10;
      13'h1e42: color = 2'b10;
      13'h1e43: color = 2'b10;
      13'h1e44: color = 2'b10;
      13'h1e45: color = 2'b10;
      13'h1e46: color = 2'b10;
      13'h1e47: color = 2'b10;
      13'h1e48: color = 2'b10;
      13'h1e49: color = 2'b10;
      13'h1e4a: color = 2'b10;
      13'h1e4b: color = 2'b10;
      13'h1e4c: color = 2'b10;
      13'h1e4d: color = 2'b10;
      13'h1e4e: color = 2'b10;
      13'h1e4f: color = 2'b10;
      13'h1e50: color = 2'b10;
      13'h1e51: color = 2'b10;
      13'h1e52: color = 2'b10;
      13'h1e53: color = 2'b10;
      13'h1e54: color = 2'b00;
      13'h1e55: color = 2'b00;
      13'h1e56: color = 2'b00;
      13'h1e57: color = 2'b00;
      13'h1e58: color = 2'b00;
      13'h1e59: color = 2'b00;
      13'h1e5a: color = 2'b00;
      13'h1e5b: color = 2'b00;
      13'h1e5c: color = 2'b00;
      13'h1e5d: color = 2'b00;
      13'h1e5e: color = 2'b11;
      13'h1e5f: color = 2'b11;
      13'h1e60: color = 2'b11;
      13'h1e61: color = 2'b11;
      13'h1e62: color = 2'b11;
      13'h1e63: color = 2'b11;
      13'h1e64: color = 2'b00;
      13'h1e65: color = 2'b00;
      13'h1e66: color = 2'b10;
      13'h1e67: color = 2'b10;
      13'h1e68: color = 2'b00;
      13'h1e69: color = 2'b00;
      13'h1e6a: color = 2'b11;
      13'h1e6b: color = 2'b11;
      13'h1e6c: color = 2'b11;
      13'h1e6d: color = 2'b11;
      13'h1e6e: color = 2'b11;
      13'h1e6f: color = 2'b11;
      13'h1e70: color = 2'b11;
      13'h1e71: color = 2'b11;
      13'h1e72: color = 2'b11;
      13'h1e73: color = 2'b11;
      13'h1e74: color = 2'b10;
      13'h1e75: color = 2'b10;
      13'h1e76: color = 2'b00;
      13'h1e77: color = 2'b00;
      13'h1e78: color = 2'b10;
      13'h1e79: color = 2'b10;
      13'h1e7a: color = 2'b00;
      13'h1e7b: color = 2'b00;
      13'h1e7c: color = 2'b11;
      13'h1e7d: color = 2'b11;
      13'h1e7e: color = 2'b11;
      13'h1e7f: color = 2'b11;
      13'h1e80: color = 2'b11;
      13'h1e81: color = 2'b11;
      13'h1e82: color = 2'b11;
      13'h1e83: color = 2'b11;
      13'h1e84: color = 2'b00;
      13'h1e85: color = 2'b00;
      13'h1e86: color = 2'b10;
      13'h1e87: color = 2'b10;
      13'h1e88: color = 2'b00;
      13'h1e89: color = 2'b00;
      13'h1e8a: color = 2'b11;
      13'h1e8b: color = 2'b11;
      13'h1e8c: color = 2'b11;
      13'h1e8d: color = 2'b11;
      13'h1e8e: color = 2'b11;
      13'h1e8f: color = 2'b11;
      13'h1e90: color = 2'b11;
      13'h1e91: color = 2'b11;
      13'h1e92: color = 2'b11;
      13'h1e93: color = 2'b11;
      13'h1e94: color = 2'b10;
      13'h1e95: color = 2'b10;
      13'h1e96: color = 2'b00;
      13'h1e97: color = 2'b00;
      13'h1e98: color = 2'b10;
      13'h1e99: color = 2'b10;
      13'h1e9a: color = 2'b00;
      13'h1e9b: color = 2'b00;
      13'h1e9c: color = 2'b11;
      13'h1e9d: color = 2'b11;
      13'h1e9e: color = 2'b11;
      13'h1e9f: color = 2'b11;
      13'h1ea0: color = 2'b11;
      13'h1ea1: color = 2'b11;
      13'h1ea2: color = 2'b00;
      13'h1ea3: color = 2'b00;
      13'h1ea4: color = 2'b00;
      13'h1ea5: color = 2'b00;
      13'h1ea6: color = 2'b00;
      13'h1ea7: color = 2'b00;
      13'h1ea8: color = 2'b00;
      13'h1ea9: color = 2'b00;
      13'h1eaa: color = 2'b00;
      13'h1eab: color = 2'b00;
      13'h1eac: color = 2'b10;
      13'h1ead: color = 2'b10;
      13'h1eae: color = 2'b10;
      13'h1eaf: color = 2'b10;
      13'h1eb0: color = 2'b10;
      13'h1eb1: color = 2'b10;
      13'h1eb2: color = 2'b10;
      13'h1eb3: color = 2'b10;
      13'h1eb4: color = 2'b10;
      13'h1eb5: color = 2'b10;
      13'h1eb6: color = 2'b10;
      13'h1eb7: color = 2'b10;
      13'h1eb8: color = 2'b10;
      13'h1eb9: color = 2'b10;
      13'h1eba: color = 2'b10;
      13'h1ebb: color = 2'b10;
      13'h1ebc: color = 2'b10;
      13'h1ebd: color = 2'b10;
      13'h1ebe: color = 2'b10;
      13'h1ebf: color = 2'b10;
      13'h1ec0: color = 2'b10;
      13'h1ec1: color = 2'b10;
      13'h1ec2: color = 2'b10;
      13'h1ec3: color = 2'b10;
      13'h1ec4: color = 2'b10;
      13'h1ec5: color = 2'b10;
      13'h1ec6: color = 2'b10;
      13'h1ec7: color = 2'b10;
      13'h1ec8: color = 2'b10;
      13'h1ec9: color = 2'b10;
      13'h1eca: color = 2'b10;
      13'h1ecb: color = 2'b10;
      13'h1ecc: color = 2'b10;
      13'h1ecd: color = 2'b10;
      13'h1ece: color = 2'b10;
      13'h1ecf: color = 2'b10;
      13'h1ed0: color = 2'b10;
      13'h1ed1: color = 2'b10;
      13'h1ed2: color = 2'b10;
      13'h1ed3: color = 2'b10;
      13'h1ed4: color = 2'b00;
      13'h1ed5: color = 2'b00;
      13'h1ed6: color = 2'b00;
      13'h1ed7: color = 2'b00;
      13'h1ed8: color = 2'b00;
      13'h1ed9: color = 2'b00;
      13'h1eda: color = 2'b00;
      13'h1edb: color = 2'b00;
      13'h1edc: color = 2'b00;
      13'h1edd: color = 2'b00;
      13'h1ede: color = 2'b11;
      13'h1edf: color = 2'b11;
      13'h1ee0: color = 2'b11;
      13'h1ee1: color = 2'b11;
      13'h1ee2: color = 2'b11;
      13'h1ee3: color = 2'b11;
      13'h1ee4: color = 2'b00;
      13'h1ee5: color = 2'b00;
      13'h1ee6: color = 2'b10;
      13'h1ee7: color = 2'b10;
      13'h1ee8: color = 2'b00;
      13'h1ee9: color = 2'b00;
      13'h1eea: color = 2'b11;
      13'h1eeb: color = 2'b11;
      13'h1eec: color = 2'b11;
      13'h1eed: color = 2'b11;
      13'h1eee: color = 2'b11;
      13'h1eef: color = 2'b11;
      13'h1ef0: color = 2'b11;
      13'h1ef1: color = 2'b11;
      13'h1ef2: color = 2'b11;
      13'h1ef3: color = 2'b11;
      13'h1ef4: color = 2'b10;
      13'h1ef5: color = 2'b10;
      13'h1ef6: color = 2'b00;
      13'h1ef7: color = 2'b00;
      13'h1ef8: color = 2'b10;
      13'h1ef9: color = 2'b10;
      13'h1efa: color = 2'b00;
      13'h1efb: color = 2'b00;
      13'h1efc: color = 2'b11;
      13'h1efd: color = 2'b11;
      13'h1efe: color = 2'b11;
      13'h1eff: color = 2'b11;
      13'h1f00: color = 2'b11;
      13'h1f01: color = 2'b11;
      13'h1f02: color = 2'b11;
      13'h1f03: color = 2'b11;
      13'h1f04: color = 2'b00;
      13'h1f05: color = 2'b00;
      13'h1f06: color = 2'b00;
      13'h1f07: color = 2'b00;
      13'h1f08: color = 2'b00;
      13'h1f09: color = 2'b00;
      13'h1f0a: color = 2'b11;
      13'h1f0b: color = 2'b11;
      13'h1f0c: color = 2'b11;
      13'h1f0d: color = 2'b11;
      13'h1f0e: color = 2'b11;
      13'h1f0f: color = 2'b11;
      13'h1f10: color = 2'b11;
      13'h1f11: color = 2'b11;
      13'h1f12: color = 2'b11;
      13'h1f13: color = 2'b11;
      13'h1f14: color = 2'b11;
      13'h1f15: color = 2'b11;
      13'h1f16: color = 2'b00;
      13'h1f17: color = 2'b00;
      13'h1f18: color = 2'b00;
      13'h1f19: color = 2'b00;
      13'h1f1a: color = 2'b00;
      13'h1f1b: color = 2'b00;
      13'h1f1c: color = 2'b11;
      13'h1f1d: color = 2'b11;
      13'h1f1e: color = 2'b11;
      13'h1f1f: color = 2'b11;
      13'h1f20: color = 2'b11;
      13'h1f21: color = 2'b11;
      13'h1f22: color = 2'b11;
      13'h1f23: color = 2'b11;
      13'h1f24: color = 2'b11;
      13'h1f25: color = 2'b11;
      13'h1f26: color = 2'b10;
      13'h1f27: color = 2'b10;
      13'h1f28: color = 2'b11;
      13'h1f29: color = 2'b11;
      13'h1f2a: color = 2'b11;
      13'h1f2b: color = 2'b11;
      13'h1f2c: color = 2'b11;
      13'h1f2d: color = 2'b11;
      13'h1f2e: color = 2'b11;
      13'h1f2f: color = 2'b11;
      13'h1f30: color = 2'b11;
      13'h1f31: color = 2'b11;
      13'h1f32: color = 2'b11;
      13'h1f33: color = 2'b11;
      13'h1f34: color = 2'b11;
      13'h1f35: color = 2'b11;
      13'h1f36: color = 2'b10;
      13'h1f37: color = 2'b10;
      13'h1f38: color = 2'b11;
      13'h1f39: color = 2'b11;
      13'h1f3a: color = 2'b11;
      13'h1f3b: color = 2'b11;
      13'h1f3c: color = 2'b11;
      13'h1f3d: color = 2'b11;
      13'h1f3e: color = 2'b11;
      13'h1f3f: color = 2'b11;
      13'h1f40: color = 2'b11;
      13'h1f41: color = 2'b11;
      13'h1f42: color = 2'b11;
      13'h1f43: color = 2'b11;
      13'h1f44: color = 2'b11;
      13'h1f45: color = 2'b11;
      13'h1f46: color = 2'b10;
      13'h1f47: color = 2'b10;
      13'h1f48: color = 2'b11;
      13'h1f49: color = 2'b11;
      13'h1f4a: color = 2'b11;
      13'h1f4b: color = 2'b11;
      13'h1f4c: color = 2'b11;
      13'h1f4d: color = 2'b11;
      13'h1f4e: color = 2'b11;
      13'h1f4f: color = 2'b11;
      13'h1f50: color = 2'b11;
      13'h1f51: color = 2'b11;
      13'h1f52: color = 2'b11;
      13'h1f53: color = 2'b11;
      13'h1f54: color = 2'b11;
      13'h1f55: color = 2'b11;
      13'h1f56: color = 2'b10;
      13'h1f57: color = 2'b10;
      13'h1f58: color = 2'b11;
      13'h1f59: color = 2'b11;
      13'h1f5a: color = 2'b11;
      13'h1f5b: color = 2'b11;
      13'h1f5c: color = 2'b11;
      13'h1f5d: color = 2'b11;
      13'h1f5e: color = 2'b11;
      13'h1f5f: color = 2'b11;
      13'h1f60: color = 2'b11;
      13'h1f61: color = 2'b11;
      13'h1f62: color = 2'b11;
      13'h1f63: color = 2'b11;
      13'h1f64: color = 2'b00;
      13'h1f65: color = 2'b00;
      13'h1f66: color = 2'b00;
      13'h1f67: color = 2'b00;
      13'h1f68: color = 2'b00;
      13'h1f69: color = 2'b00;
      13'h1f6a: color = 2'b11;
      13'h1f6b: color = 2'b11;
      13'h1f6c: color = 2'b11;
      13'h1f6d: color = 2'b11;
      13'h1f6e: color = 2'b11;
      13'h1f6f: color = 2'b11;
      13'h1f70: color = 2'b11;
      13'h1f71: color = 2'b11;
      13'h1f72: color = 2'b11;
      13'h1f73: color = 2'b11;
      13'h1f74: color = 2'b11;
      13'h1f75: color = 2'b11;
      13'h1f76: color = 2'b00;
      13'h1f77: color = 2'b00;
      13'h1f78: color = 2'b00;
      13'h1f79: color = 2'b00;
      13'h1f7a: color = 2'b00;
      13'h1f7b: color = 2'b00;
      13'h1f7c: color = 2'b11;
      13'h1f7d: color = 2'b11;
      13'h1f7e: color = 2'b11;
      13'h1f7f: color = 2'b11;
      13'h1f80: color = 2'b11;
      13'h1f81: color = 2'b11;
      13'h1f82: color = 2'b11;
      13'h1f83: color = 2'b11;
      13'h1f84: color = 2'b00;
      13'h1f85: color = 2'b00;
      13'h1f86: color = 2'b00;
      13'h1f87: color = 2'b00;
      13'h1f88: color = 2'b00;
      13'h1f89: color = 2'b00;
      13'h1f8a: color = 2'b11;
      13'h1f8b: color = 2'b11;
      13'h1f8c: color = 2'b11;
      13'h1f8d: color = 2'b11;
      13'h1f8e: color = 2'b11;
      13'h1f8f: color = 2'b11;
      13'h1f90: color = 2'b11;
      13'h1f91: color = 2'b11;
      13'h1f92: color = 2'b11;
      13'h1f93: color = 2'b11;
      13'h1f94: color = 2'b11;
      13'h1f95: color = 2'b11;
      13'h1f96: color = 2'b00;
      13'h1f97: color = 2'b00;
      13'h1f98: color = 2'b00;
      13'h1f99: color = 2'b00;
      13'h1f9a: color = 2'b00;
      13'h1f9b: color = 2'b00;
      13'h1f9c: color = 2'b11;
      13'h1f9d: color = 2'b11;
      13'h1f9e: color = 2'b11;
      13'h1f9f: color = 2'b11;
      13'h1fa0: color = 2'b11;
      13'h1fa1: color = 2'b11;
      13'h1fa2: color = 2'b11;
      13'h1fa3: color = 2'b11;
      13'h1fa4: color = 2'b11;
      13'h1fa5: color = 2'b11;
      13'h1fa6: color = 2'b10;
      13'h1fa7: color = 2'b10;
      13'h1fa8: color = 2'b11;
      13'h1fa9: color = 2'b11;
      13'h1faa: color = 2'b11;
      13'h1fab: color = 2'b11;
      13'h1fac: color = 2'b11;
      13'h1fad: color = 2'b11;
      13'h1fae: color = 2'b11;
      13'h1faf: color = 2'b11;
      13'h1fb0: color = 2'b11;
      13'h1fb1: color = 2'b11;
      13'h1fb2: color = 2'b11;
      13'h1fb3: color = 2'b11;
      13'h1fb4: color = 2'b11;
      13'h1fb5: color = 2'b11;
      13'h1fb6: color = 2'b10;
      13'h1fb7: color = 2'b10;
      13'h1fb8: color = 2'b11;
      13'h1fb9: color = 2'b11;
      13'h1fba: color = 2'b11;
      13'h1fbb: color = 2'b11;
      13'h1fbc: color = 2'b11;
      13'h1fbd: color = 2'b11;
      13'h1fbe: color = 2'b11;
      13'h1fbf: color = 2'b11;
      13'h1fc0: color = 2'b11;
      13'h1fc1: color = 2'b11;
      13'h1fc2: color = 2'b11;
      13'h1fc3: color = 2'b11;
      13'h1fc4: color = 2'b11;
      13'h1fc5: color = 2'b11;
      13'h1fc6: color = 2'b10;
      13'h1fc7: color = 2'b10;
      13'h1fc8: color = 2'b11;
      13'h1fc9: color = 2'b11;
      13'h1fca: color = 2'b11;
      13'h1fcb: color = 2'b11;
      13'h1fcc: color = 2'b11;
      13'h1fcd: color = 2'b11;
      13'h1fce: color = 2'b11;
      13'h1fcf: color = 2'b11;
      13'h1fd0: color = 2'b11;
      13'h1fd1: color = 2'b11;
      13'h1fd2: color = 2'b11;
      13'h1fd3: color = 2'b11;
      13'h1fd4: color = 2'b11;
      13'h1fd5: color = 2'b11;
      13'h1fd6: color = 2'b10;
      13'h1fd7: color = 2'b10;
      13'h1fd8: color = 2'b11;
      13'h1fd9: color = 2'b11;
      13'h1fda: color = 2'b11;
      13'h1fdb: color = 2'b11;
      13'h1fdc: color = 2'b11;
      13'h1fdd: color = 2'b11;
      13'h1fde: color = 2'b11;
      13'h1fdf: color = 2'b11;
      13'h1fe0: color = 2'b11;
      13'h1fe1: color = 2'b11;
      13'h1fe2: color = 2'b11;
      13'h1fe3: color = 2'b11;
      13'h1fe4: color = 2'b00;
      13'h1fe5: color = 2'b00;
      13'h1fe6: color = 2'b00;
      13'h1fe7: color = 2'b00;
      13'h1fe8: color = 2'b00;
      13'h1fe9: color = 2'b00;
      13'h1fea: color = 2'b11;
      13'h1feb: color = 2'b11;
      13'h1fec: color = 2'b11;
      13'h1fed: color = 2'b11;
      13'h1fee: color = 2'b11;
      13'h1fef: color = 2'b11;
      13'h1ff0: color = 2'b11;
      13'h1ff1: color = 2'b11;
      13'h1ff2: color = 2'b11;
      13'h1ff3: color = 2'b11;
      13'h1ff4: color = 2'b11;
      13'h1ff5: color = 2'b11;
      13'h1ff6: color = 2'b00;
      13'h1ff7: color = 2'b00;
      13'h1ff8: color = 2'b00;
      13'h1ff9: color = 2'b00;
      13'h1ffa: color = 2'b00;
      13'h1ffb: color = 2'b00;
      13'h1ffc: color = 2'b11;
      13'h1ffd: color = 2'b11;
      13'h1ffe: color = 2'b11;
      13'h1fff: color = 2'b11;
   endcase
end
endmodule
