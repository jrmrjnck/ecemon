
`define UP_ARROW    8'h75
`define DOWN_ARROW  8'h72
`define RIGHT_ARROW 8'h74
`define LEFT_ARROW  8'h6B
`define ENTER       8'h5A
`define KEY_A       8'h1C
`define KEY_B       8'h32

`define BLACK 2'b00
`define DARK  2'b01
`define LIGHT 2'b10
`define WHITE 2'b11

`define SPLASH_STATE 3'd0
`define INTRO_STATE  3'd1
`define CEL_STATE    3'd2
`define COMP_STATE   3'd3
`define ATTACK_STATE  3'd4
`define QUESTION_STATE 3'd5

`define PROF_TOM 3'd0
`define PROF_JASON 3'd1
`define PROF_PAUL 3'd2
`define PROF_MARK 3'd3
