module Paul
(
   input            clock, 
   input      [7:0] x,
   input      [7:0] y, 
   input      [7:0] loc_x, 
   input      [7:0] loc_y, 
   output reg       on,
   output reg [1:0] color
);

   localparam WIDTH = 8'd128,
              HEIGHT = 8'd128;

   // Buffer the scan coordinates to synchronize
   // with the ROM data output
   always @( posedge clock ) begin
    on <= (x >= loc_x && x <= (loc_x+(WIDTH-1)))
          && (y >= loc_y && y <= (loc_y+(HEIGHT-1)));
   end

   reg [13:0] addr;
   always @( posedge clock )
      addr <= {y[6:0]-loc_y[6:0],x[6:0]-loc_x[6:0]};
   
always @(*) begin
	case( addr )
		14'h0000: color = 2'b11;
		14'h0001: color = 2'b11;
		14'h0002: color = 2'b11;
		14'h0003: color = 2'b11;
		14'h0004: color = 2'b11;
		14'h0005: color = 2'b11;
		14'h0006: color = 2'b11;
		14'h0007: color = 2'b11;
		14'h0008: color = 2'b11;
		14'h0009: color = 2'b11;
		14'h000a: color = 2'b11;
		14'h000b: color = 2'b11;
		14'h000c: color = 2'b11;
		14'h000d: color = 2'b11;
		14'h000e: color = 2'b11;
		14'h000f: color = 2'b11;
		14'h0010: color = 2'b11;
		14'h0011: color = 2'b11;
		14'h0012: color = 2'b11;
		14'h0013: color = 2'b11;
		14'h0014: color = 2'b11;
		14'h0015: color = 2'b11;
		14'h0016: color = 2'b11;
		14'h0017: color = 2'b11;
		14'h0018: color = 2'b11;
		14'h0019: color = 2'b11;
		14'h001a: color = 2'b11;
		14'h001b: color = 2'b11;
		14'h001c: color = 2'b11;
		14'h001d: color = 2'b11;
		14'h001e: color = 2'b11;
		14'h001f: color = 2'b11;
		14'h0020: color = 2'b11;
		14'h0021: color = 2'b11;
		14'h0022: color = 2'b11;
		14'h0023: color = 2'b11;
		14'h0024: color = 2'b11;
		14'h0025: color = 2'b11;
		14'h0026: color = 2'b11;
		14'h0027: color = 2'b11;
		14'h0028: color = 2'b11;
		14'h0029: color = 2'b11;
		14'h002a: color = 2'b11;
		14'h002b: color = 2'b11;
		14'h002c: color = 2'b11;
		14'h002d: color = 2'b11;
		14'h002e: color = 2'b11;
		14'h002f: color = 2'b11;
		14'h0030: color = 2'b11;
		14'h0031: color = 2'b11;
		14'h0032: color = 2'b11;
		14'h0033: color = 2'b11;
		14'h0034: color = 2'b11;
		14'h0035: color = 2'b11;
		14'h0036: color = 2'b11;
		14'h0037: color = 2'b11;
		14'h0038: color = 2'b11;
		14'h0039: color = 2'b11;
		14'h003a: color = 2'b11;
		14'h003b: color = 2'b11;
		14'h003c: color = 2'b11;
		14'h003d: color = 2'b11;
		14'h003e: color = 2'b11;
		14'h003f: color = 2'b11;
		14'h0040: color = 2'b11;
		14'h0041: color = 2'b11;
		14'h0042: color = 2'b11;
		14'h0043: color = 2'b11;
		14'h0044: color = 2'b11;
		14'h0045: color = 2'b11;
		14'h0046: color = 2'b11;
		14'h0047: color = 2'b11;
		14'h0048: color = 2'b11;
		14'h0049: color = 2'b11;
		14'h004a: color = 2'b11;
		14'h004b: color = 2'b11;
		14'h004c: color = 2'b11;
		14'h004d: color = 2'b11;
		14'h004e: color = 2'b11;
		14'h004f: color = 2'b11;
		14'h0050: color = 2'b11;
		14'h0051: color = 2'b11;
		14'h0052: color = 2'b11;
		14'h0053: color = 2'b11;
		14'h0054: color = 2'b11;
		14'h0055: color = 2'b11;
		14'h0056: color = 2'b11;
		14'h0057: color = 2'b11;
		14'h0058: color = 2'b11;
		14'h0059: color = 2'b11;
		14'h005a: color = 2'b11;
		14'h005b: color = 2'b11;
		14'h005c: color = 2'b11;
		14'h005d: color = 2'b11;
		14'h005e: color = 2'b11;
		14'h005f: color = 2'b11;
		14'h0060: color = 2'b11;
		14'h0061: color = 2'b11;
		14'h0062: color = 2'b11;
		14'h0063: color = 2'b11;
		14'h0064: color = 2'b11;
		14'h0065: color = 2'b11;
		14'h0066: color = 2'b11;
		14'h0067: color = 2'b11;
		14'h0068: color = 2'b11;
		14'h0069: color = 2'b11;
		14'h006a: color = 2'b11;
		14'h006b: color = 2'b11;
		14'h006c: color = 2'b11;
		14'h006d: color = 2'b11;
		14'h006e: color = 2'b11;
		14'h006f: color = 2'b11;
		14'h0070: color = 2'b11;
		14'h0071: color = 2'b11;
		14'h0072: color = 2'b11;
		14'h0073: color = 2'b11;
		14'h0074: color = 2'b11;
		14'h0075: color = 2'b11;
		14'h0076: color = 2'b11;
		14'h0077: color = 2'b11;
		14'h0078: color = 2'b11;
		14'h0079: color = 2'b11;
		14'h007a: color = 2'b11;
		14'h007b: color = 2'b11;
		14'h007c: color = 2'b11;
		14'h007d: color = 2'b11;
		14'h007e: color = 2'b11;
		14'h007f: color = 2'b11;
		14'h0080: color = 2'b11;
		14'h0081: color = 2'b11;
		14'h0082: color = 2'b11;
		14'h0083: color = 2'b11;
		14'h0084: color = 2'b11;
		14'h0085: color = 2'b11;
		14'h0086: color = 2'b11;
		14'h0087: color = 2'b11;
		14'h0088: color = 2'b11;
		14'h0089: color = 2'b11;
		14'h008a: color = 2'b11;
		14'h008b: color = 2'b11;
		14'h008c: color = 2'b11;
		14'h008d: color = 2'b11;
		14'h008e: color = 2'b11;
		14'h008f: color = 2'b11;
		14'h0090: color = 2'b11;
		14'h0091: color = 2'b11;
		14'h0092: color = 2'b11;
		14'h0093: color = 2'b11;
		14'h0094: color = 2'b11;
		14'h0095: color = 2'b11;
		14'h0096: color = 2'b11;
		14'h0097: color = 2'b11;
		14'h0098: color = 2'b11;
		14'h0099: color = 2'b11;
		14'h009a: color = 2'b11;
		14'h009b: color = 2'b11;
		14'h009c: color = 2'b11;
		14'h009d: color = 2'b11;
		14'h009e: color = 2'b11;
		14'h009f: color = 2'b11;
		14'h00a0: color = 2'b11;
		14'h00a1: color = 2'b11;
		14'h00a2: color = 2'b11;
		14'h00a3: color = 2'b11;
		14'h00a4: color = 2'b11;
		14'h00a5: color = 2'b11;
		14'h00a6: color = 2'b11;
		14'h00a7: color = 2'b11;
		14'h00a8: color = 2'b11;
		14'h00a9: color = 2'b11;
		14'h00aa: color = 2'b11;
		14'h00ab: color = 2'b11;
		14'h00ac: color = 2'b11;
		14'h00ad: color = 2'b11;
		14'h00ae: color = 2'b11;
		14'h00af: color = 2'b11;
		14'h00b0: color = 2'b11;
		14'h00b1: color = 2'b11;
		14'h00b2: color = 2'b11;
		14'h00b3: color = 2'b11;
		14'h00b4: color = 2'b11;
		14'h00b5: color = 2'b11;
		14'h00b6: color = 2'b11;
		14'h00b7: color = 2'b11;
		14'h00b8: color = 2'b11;
		14'h00b9: color = 2'b11;
		14'h00ba: color = 2'b11;
		14'h00bb: color = 2'b11;
		14'h00bc: color = 2'b11;
		14'h00bd: color = 2'b11;
		14'h00be: color = 2'b11;
		14'h00bf: color = 2'b11;
		14'h00c0: color = 2'b11;
		14'h00c1: color = 2'b11;
		14'h00c2: color = 2'b11;
		14'h00c3: color = 2'b11;
		14'h00c4: color = 2'b11;
		14'h00c5: color = 2'b11;
		14'h00c6: color = 2'b11;
		14'h00c7: color = 2'b11;
		14'h00c8: color = 2'b11;
		14'h00c9: color = 2'b11;
		14'h00ca: color = 2'b11;
		14'h00cb: color = 2'b11;
		14'h00cc: color = 2'b11;
		14'h00cd: color = 2'b11;
		14'h00ce: color = 2'b11;
		14'h00cf: color = 2'b11;
		14'h00d0: color = 2'b11;
		14'h00d1: color = 2'b11;
		14'h00d2: color = 2'b11;
		14'h00d3: color = 2'b11;
		14'h00d4: color = 2'b11;
		14'h00d5: color = 2'b11;
		14'h00d6: color = 2'b11;
		14'h00d7: color = 2'b11;
		14'h00d8: color = 2'b11;
		14'h00d9: color = 2'b11;
		14'h00da: color = 2'b11;
		14'h00db: color = 2'b11;
		14'h00dc: color = 2'b11;
		14'h00dd: color = 2'b11;
		14'h00de: color = 2'b11;
		14'h00df: color = 2'b11;
		14'h00e0: color = 2'b11;
		14'h00e1: color = 2'b11;
		14'h00e2: color = 2'b11;
		14'h00e3: color = 2'b11;
		14'h00e4: color = 2'b11;
		14'h00e5: color = 2'b11;
		14'h00e6: color = 2'b11;
		14'h00e7: color = 2'b11;
		14'h00e8: color = 2'b11;
		14'h00e9: color = 2'b11;
		14'h00ea: color = 2'b11;
		14'h00eb: color = 2'b11;
		14'h00ec: color = 2'b11;
		14'h00ed: color = 2'b11;
		14'h00ee: color = 2'b11;
		14'h00ef: color = 2'b11;
		14'h00f0: color = 2'b11;
		14'h00f1: color = 2'b11;
		14'h00f2: color = 2'b11;
		14'h00f3: color = 2'b11;
		14'h00f4: color = 2'b11;
		14'h00f5: color = 2'b11;
		14'h00f6: color = 2'b11;
		14'h00f7: color = 2'b11;
		14'h00f8: color = 2'b11;
		14'h00f9: color = 2'b11;
		14'h00fa: color = 2'b11;
		14'h00fb: color = 2'b11;
		14'h00fc: color = 2'b11;
		14'h00fd: color = 2'b11;
		14'h00fe: color = 2'b11;
		14'h00ff: color = 2'b11;
		14'h0100: color = 2'b11;
		14'h0101: color = 2'b11;
		14'h0102: color = 2'b11;
		14'h0103: color = 2'b11;
		14'h0104: color = 2'b11;
		14'h0105: color = 2'b11;
		14'h0106: color = 2'b11;
		14'h0107: color = 2'b11;
		14'h0108: color = 2'b11;
		14'h0109: color = 2'b11;
		14'h010a: color = 2'b11;
		14'h010b: color = 2'b11;
		14'h010c: color = 2'b11;
		14'h010d: color = 2'b11;
		14'h010e: color = 2'b11;
		14'h010f: color = 2'b11;
		14'h0110: color = 2'b11;
		14'h0111: color = 2'b11;
		14'h0112: color = 2'b11;
		14'h0113: color = 2'b11;
		14'h0114: color = 2'b11;
		14'h0115: color = 2'b11;
		14'h0116: color = 2'b11;
		14'h0117: color = 2'b11;
		14'h0118: color = 2'b11;
		14'h0119: color = 2'b11;
		14'h011a: color = 2'b11;
		14'h011b: color = 2'b11;
		14'h011c: color = 2'b11;
		14'h011d: color = 2'b11;
		14'h011e: color = 2'b11;
		14'h011f: color = 2'b11;
		14'h0120: color = 2'b11;
		14'h0121: color = 2'b11;
		14'h0122: color = 2'b11;
		14'h0123: color = 2'b11;
		14'h0124: color = 2'b11;
		14'h0125: color = 2'b11;
		14'h0126: color = 2'b11;
		14'h0127: color = 2'b11;
		14'h0128: color = 2'b11;
		14'h0129: color = 2'b11;
		14'h012a: color = 2'b11;
		14'h012b: color = 2'b11;
		14'h012c: color = 2'b11;
		14'h012d: color = 2'b11;
		14'h012e: color = 2'b11;
		14'h012f: color = 2'b11;
		14'h0130: color = 2'b11;
		14'h0131: color = 2'b11;
		14'h0132: color = 2'b11;
		14'h0133: color = 2'b11;
		14'h0134: color = 2'b11;
		14'h0135: color = 2'b11;
		14'h0136: color = 2'b11;
		14'h0137: color = 2'b11;
		14'h0138: color = 2'b11;
		14'h0139: color = 2'b11;
		14'h013a: color = 2'b11;
		14'h013b: color = 2'b11;
		14'h013c: color = 2'b11;
		14'h013d: color = 2'b11;
		14'h013e: color = 2'b11;
		14'h013f: color = 2'b11;
		14'h0140: color = 2'b11;
		14'h0141: color = 2'b11;
		14'h0142: color = 2'b11;
		14'h0143: color = 2'b11;
		14'h0144: color = 2'b11;
		14'h0145: color = 2'b11;
		14'h0146: color = 2'b11;
		14'h0147: color = 2'b11;
		14'h0148: color = 2'b11;
		14'h0149: color = 2'b11;
		14'h014a: color = 2'b11;
		14'h014b: color = 2'b11;
		14'h014c: color = 2'b11;
		14'h014d: color = 2'b11;
		14'h014e: color = 2'b11;
		14'h014f: color = 2'b11;
		14'h0150: color = 2'b11;
		14'h0151: color = 2'b11;
		14'h0152: color = 2'b11;
		14'h0153: color = 2'b11;
		14'h0154: color = 2'b11;
		14'h0155: color = 2'b11;
		14'h0156: color = 2'b11;
		14'h0157: color = 2'b11;
		14'h0158: color = 2'b11;
		14'h0159: color = 2'b11;
		14'h015a: color = 2'b11;
		14'h015b: color = 2'b11;
		14'h015c: color = 2'b11;
		14'h015d: color = 2'b11;
		14'h015e: color = 2'b11;
		14'h015f: color = 2'b11;
		14'h0160: color = 2'b11;
		14'h0161: color = 2'b11;
		14'h0162: color = 2'b11;
		14'h0163: color = 2'b11;
		14'h0164: color = 2'b11;
		14'h0165: color = 2'b11;
		14'h0166: color = 2'b11;
		14'h0167: color = 2'b11;
		14'h0168: color = 2'b11;
		14'h0169: color = 2'b11;
		14'h016a: color = 2'b11;
		14'h016b: color = 2'b11;
		14'h016c: color = 2'b11;
		14'h016d: color = 2'b11;
		14'h016e: color = 2'b11;
		14'h016f: color = 2'b11;
		14'h0170: color = 2'b11;
		14'h0171: color = 2'b11;
		14'h0172: color = 2'b11;
		14'h0173: color = 2'b11;
		14'h0174: color = 2'b11;
		14'h0175: color = 2'b11;
		14'h0176: color = 2'b11;
		14'h0177: color = 2'b11;
		14'h0178: color = 2'b11;
		14'h0179: color = 2'b11;
		14'h017a: color = 2'b11;
		14'h017b: color = 2'b11;
		14'h017c: color = 2'b11;
		14'h017d: color = 2'b11;
		14'h017e: color = 2'b11;
		14'h017f: color = 2'b11;
		14'h0180: color = 2'b11;
		14'h0181: color = 2'b11;
		14'h0182: color = 2'b11;
		14'h0183: color = 2'b11;
		14'h0184: color = 2'b11;
		14'h0185: color = 2'b11;
		14'h0186: color = 2'b11;
		14'h0187: color = 2'b11;
		14'h0188: color = 2'b11;
		14'h0189: color = 2'b11;
		14'h018a: color = 2'b11;
		14'h018b: color = 2'b11;
		14'h018c: color = 2'b11;
		14'h018d: color = 2'b11;
		14'h018e: color = 2'b11;
		14'h018f: color = 2'b11;
		14'h0190: color = 2'b11;
		14'h0191: color = 2'b11;
		14'h0192: color = 2'b11;
		14'h0193: color = 2'b11;
		14'h0194: color = 2'b11;
		14'h0195: color = 2'b11;
		14'h0196: color = 2'b11;
		14'h0197: color = 2'b11;
		14'h0198: color = 2'b11;
		14'h0199: color = 2'b11;
		14'h019a: color = 2'b11;
		14'h019b: color = 2'b11;
		14'h019c: color = 2'b11;
		14'h019d: color = 2'b11;
		14'h019e: color = 2'b11;
		14'h019f: color = 2'b11;
		14'h01a0: color = 2'b11;
		14'h01a1: color = 2'b11;
		14'h01a2: color = 2'b11;
		14'h01a3: color = 2'b11;
		14'h01a4: color = 2'b11;
		14'h01a5: color = 2'b11;
		14'h01a6: color = 2'b11;
		14'h01a7: color = 2'b11;
		14'h01a8: color = 2'b11;
		14'h01a9: color = 2'b11;
		14'h01aa: color = 2'b11;
		14'h01ab: color = 2'b11;
		14'h01ac: color = 2'b11;
		14'h01ad: color = 2'b11;
		14'h01ae: color = 2'b11;
		14'h01af: color = 2'b11;
		14'h01b0: color = 2'b11;
		14'h01b1: color = 2'b11;
		14'h01b2: color = 2'b11;
		14'h01b3: color = 2'b11;
		14'h01b4: color = 2'b11;
		14'h01b5: color = 2'b11;
		14'h01b6: color = 2'b11;
		14'h01b7: color = 2'b11;
		14'h01b8: color = 2'b11;
		14'h01b9: color = 2'b11;
		14'h01ba: color = 2'b11;
		14'h01bb: color = 2'b11;
		14'h01bc: color = 2'b11;
		14'h01bd: color = 2'b11;
		14'h01be: color = 2'b11;
		14'h01bf: color = 2'b11;
		14'h01c0: color = 2'b11;
		14'h01c1: color = 2'b11;
		14'h01c2: color = 2'b11;
		14'h01c3: color = 2'b11;
		14'h01c4: color = 2'b11;
		14'h01c5: color = 2'b11;
		14'h01c6: color = 2'b11;
		14'h01c7: color = 2'b11;
		14'h01c8: color = 2'b11;
		14'h01c9: color = 2'b11;
		14'h01ca: color = 2'b11;
		14'h01cb: color = 2'b11;
		14'h01cc: color = 2'b11;
		14'h01cd: color = 2'b11;
		14'h01ce: color = 2'b11;
		14'h01cf: color = 2'b11;
		14'h01d0: color = 2'b11;
		14'h01d1: color = 2'b11;
		14'h01d2: color = 2'b11;
		14'h01d3: color = 2'b11;
		14'h01d4: color = 2'b11;
		14'h01d5: color = 2'b11;
		14'h01d6: color = 2'b11;
		14'h01d7: color = 2'b11;
		14'h01d8: color = 2'b11;
		14'h01d9: color = 2'b11;
		14'h01da: color = 2'b11;
		14'h01db: color = 2'b11;
		14'h01dc: color = 2'b11;
		14'h01dd: color = 2'b11;
		14'h01de: color = 2'b11;
		14'h01df: color = 2'b11;
		14'h01e0: color = 2'b11;
		14'h01e1: color = 2'b11;
		14'h01e2: color = 2'b11;
		14'h01e3: color = 2'b11;
		14'h01e4: color = 2'b11;
		14'h01e5: color = 2'b11;
		14'h01e6: color = 2'b11;
		14'h01e7: color = 2'b11;
		14'h01e8: color = 2'b11;
		14'h01e9: color = 2'b11;
		14'h01ea: color = 2'b11;
		14'h01eb: color = 2'b11;
		14'h01ec: color = 2'b11;
		14'h01ed: color = 2'b11;
		14'h01ee: color = 2'b11;
		14'h01ef: color = 2'b11;
		14'h01f0: color = 2'b11;
		14'h01f1: color = 2'b11;
		14'h01f2: color = 2'b11;
		14'h01f3: color = 2'b11;
		14'h01f4: color = 2'b11;
		14'h01f5: color = 2'b11;
		14'h01f6: color = 2'b11;
		14'h01f7: color = 2'b11;
		14'h01f8: color = 2'b11;
		14'h01f9: color = 2'b11;
		14'h01fa: color = 2'b11;
		14'h01fb: color = 2'b11;
		14'h01fc: color = 2'b11;
		14'h01fd: color = 2'b11;
		14'h01fe: color = 2'b11;
		14'h01ff: color = 2'b11;
		14'h0200: color = 2'b11;
		14'h0201: color = 2'b11;
		14'h0202: color = 2'b11;
		14'h0203: color = 2'b11;
		14'h0204: color = 2'b11;
		14'h0205: color = 2'b11;
		14'h0206: color = 2'b11;
		14'h0207: color = 2'b11;
		14'h0208: color = 2'b11;
		14'h0209: color = 2'b11;
		14'h020a: color = 2'b11;
		14'h020b: color = 2'b11;
		14'h020c: color = 2'b11;
		14'h020d: color = 2'b11;
		14'h020e: color = 2'b11;
		14'h020f: color = 2'b11;
		14'h0210: color = 2'b11;
		14'h0211: color = 2'b11;
		14'h0212: color = 2'b11;
		14'h0213: color = 2'b11;
		14'h0214: color = 2'b11;
		14'h0215: color = 2'b11;
		14'h0216: color = 2'b11;
		14'h0217: color = 2'b11;
		14'h0218: color = 2'b11;
		14'h0219: color = 2'b11;
		14'h021a: color = 2'b11;
		14'h021b: color = 2'b11;
		14'h021c: color = 2'b11;
		14'h021d: color = 2'b11;
		14'h021e: color = 2'b11;
		14'h021f: color = 2'b11;
		14'h0220: color = 2'b11;
		14'h0221: color = 2'b11;
		14'h0222: color = 2'b11;
		14'h0223: color = 2'b11;
		14'h0224: color = 2'b11;
		14'h0225: color = 2'b11;
		14'h0226: color = 2'b11;
		14'h0227: color = 2'b11;
		14'h0228: color = 2'b11;
		14'h0229: color = 2'b11;
		14'h022a: color = 2'b11;
		14'h022b: color = 2'b11;
		14'h022c: color = 2'b11;
		14'h022d: color = 2'b11;
		14'h022e: color = 2'b11;
		14'h022f: color = 2'b11;
		14'h0230: color = 2'b11;
		14'h0231: color = 2'b11;
		14'h0232: color = 2'b11;
		14'h0233: color = 2'b11;
		14'h0234: color = 2'b11;
		14'h0235: color = 2'b11;
		14'h0236: color = 2'b11;
		14'h0237: color = 2'b11;
		14'h0238: color = 2'b11;
		14'h0239: color = 2'b11;
		14'h023a: color = 2'b11;
		14'h023b: color = 2'b11;
		14'h023c: color = 2'b11;
		14'h023d: color = 2'b11;
		14'h023e: color = 2'b11;
		14'h023f: color = 2'b11;
		14'h0240: color = 2'b11;
		14'h0241: color = 2'b11;
		14'h0242: color = 2'b11;
		14'h0243: color = 2'b11;
		14'h0244: color = 2'b11;
		14'h0245: color = 2'b10;
		14'h0246: color = 2'b01;
		14'h0247: color = 2'b10;
		14'h0248: color = 2'b10;
		14'h0249: color = 2'b10;
		14'h024a: color = 2'b10;
		14'h024b: color = 2'b11;
		14'h024c: color = 2'b10;
		14'h024d: color = 2'b11;
		14'h024e: color = 2'b11;
		14'h024f: color = 2'b11;
		14'h0250: color = 2'b11;
		14'h0251: color = 2'b11;
		14'h0252: color = 2'b11;
		14'h0253: color = 2'b11;
		14'h0254: color = 2'b11;
		14'h0255: color = 2'b11;
		14'h0256: color = 2'b11;
		14'h0257: color = 2'b11;
		14'h0258: color = 2'b11;
		14'h0259: color = 2'b11;
		14'h025a: color = 2'b11;
		14'h025b: color = 2'b11;
		14'h025c: color = 2'b11;
		14'h025d: color = 2'b11;
		14'h025e: color = 2'b11;
		14'h025f: color = 2'b11;
		14'h0260: color = 2'b11;
		14'h0261: color = 2'b11;
		14'h0262: color = 2'b11;
		14'h0263: color = 2'b11;
		14'h0264: color = 2'b11;
		14'h0265: color = 2'b11;
		14'h0266: color = 2'b11;
		14'h0267: color = 2'b11;
		14'h0268: color = 2'b11;
		14'h0269: color = 2'b11;
		14'h026a: color = 2'b11;
		14'h026b: color = 2'b11;
		14'h026c: color = 2'b11;
		14'h026d: color = 2'b11;
		14'h026e: color = 2'b11;
		14'h026f: color = 2'b11;
		14'h0270: color = 2'b11;
		14'h0271: color = 2'b11;
		14'h0272: color = 2'b11;
		14'h0273: color = 2'b11;
		14'h0274: color = 2'b11;
		14'h0275: color = 2'b11;
		14'h0276: color = 2'b11;
		14'h0277: color = 2'b11;
		14'h0278: color = 2'b11;
		14'h0279: color = 2'b11;
		14'h027a: color = 2'b11;
		14'h027b: color = 2'b11;
		14'h027c: color = 2'b11;
		14'h027d: color = 2'b11;
		14'h027e: color = 2'b11;
		14'h027f: color = 2'b11;
		14'h0280: color = 2'b11;
		14'h0281: color = 2'b11;
		14'h0282: color = 2'b11;
		14'h0283: color = 2'b11;
		14'h0284: color = 2'b11;
		14'h0285: color = 2'b11;
		14'h0286: color = 2'b11;
		14'h0287: color = 2'b11;
		14'h0288: color = 2'b11;
		14'h0289: color = 2'b11;
		14'h028a: color = 2'b11;
		14'h028b: color = 2'b11;
		14'h028c: color = 2'b11;
		14'h028d: color = 2'b11;
		14'h028e: color = 2'b11;
		14'h028f: color = 2'b11;
		14'h0290: color = 2'b11;
		14'h0291: color = 2'b11;
		14'h0292: color = 2'b11;
		14'h0293: color = 2'b11;
		14'h0294: color = 2'b11;
		14'h0295: color = 2'b11;
		14'h0296: color = 2'b11;
		14'h0297: color = 2'b11;
		14'h0298: color = 2'b11;
		14'h0299: color = 2'b11;
		14'h029a: color = 2'b11;
		14'h029b: color = 2'b11;
		14'h029c: color = 2'b11;
		14'h029d: color = 2'b11;
		14'h029e: color = 2'b11;
		14'h029f: color = 2'b11;
		14'h02a0: color = 2'b11;
		14'h02a1: color = 2'b11;
		14'h02a2: color = 2'b11;
		14'h02a3: color = 2'b11;
		14'h02a4: color = 2'b11;
		14'h02a5: color = 2'b11;
		14'h02a6: color = 2'b11;
		14'h02a7: color = 2'b11;
		14'h02a8: color = 2'b11;
		14'h02a9: color = 2'b11;
		14'h02aa: color = 2'b11;
		14'h02ab: color = 2'b11;
		14'h02ac: color = 2'b11;
		14'h02ad: color = 2'b11;
		14'h02ae: color = 2'b11;
		14'h02af: color = 2'b11;
		14'h02b0: color = 2'b11;
		14'h02b1: color = 2'b11;
		14'h02b2: color = 2'b11;
		14'h02b3: color = 2'b11;
		14'h02b4: color = 2'b11;
		14'h02b5: color = 2'b11;
		14'h02b6: color = 2'b11;
		14'h02b7: color = 2'b11;
		14'h02b8: color = 2'b11;
		14'h02b9: color = 2'b11;
		14'h02ba: color = 2'b11;
		14'h02bb: color = 2'b11;
		14'h02bc: color = 2'b11;
		14'h02bd: color = 2'b11;
		14'h02be: color = 2'b11;
		14'h02bf: color = 2'b11;
		14'h02c0: color = 2'b11;
		14'h02c1: color = 2'b01;
		14'h02c2: color = 2'b01;
		14'h02c3: color = 2'b10;
		14'h02c4: color = 2'b11;
		14'h02c5: color = 2'b00;
		14'h02c6: color = 2'b01;
		14'h02c7: color = 2'b00;
		14'h02c8: color = 2'b00;
		14'h02c9: color = 2'b00;
		14'h02ca: color = 2'b00;
		14'h02cb: color = 2'b01;
		14'h02cc: color = 2'b11;
		14'h02cd: color = 2'b00;
		14'h02ce: color = 2'b01;
		14'h02cf: color = 2'b11;
		14'h02d0: color = 2'b11;
		14'h02d1: color = 2'b11;
		14'h02d2: color = 2'b11;
		14'h02d3: color = 2'b11;
		14'h02d4: color = 2'b11;
		14'h02d5: color = 2'b11;
		14'h02d6: color = 2'b11;
		14'h02d7: color = 2'b11;
		14'h02d8: color = 2'b11;
		14'h02d9: color = 2'b11;
		14'h02da: color = 2'b11;
		14'h02db: color = 2'b11;
		14'h02dc: color = 2'b11;
		14'h02dd: color = 2'b11;
		14'h02de: color = 2'b11;
		14'h02df: color = 2'b11;
		14'h02e0: color = 2'b11;
		14'h02e1: color = 2'b11;
		14'h02e2: color = 2'b11;
		14'h02e3: color = 2'b11;
		14'h02e4: color = 2'b11;
		14'h02e5: color = 2'b11;
		14'h02e6: color = 2'b11;
		14'h02e7: color = 2'b11;
		14'h02e8: color = 2'b11;
		14'h02e9: color = 2'b11;
		14'h02ea: color = 2'b11;
		14'h02eb: color = 2'b11;
		14'h02ec: color = 2'b11;
		14'h02ed: color = 2'b11;
		14'h02ee: color = 2'b11;
		14'h02ef: color = 2'b11;
		14'h02f0: color = 2'b11;
		14'h02f1: color = 2'b11;
		14'h02f2: color = 2'b11;
		14'h02f3: color = 2'b11;
		14'h02f4: color = 2'b11;
		14'h02f5: color = 2'b11;
		14'h02f6: color = 2'b11;
		14'h02f7: color = 2'b11;
		14'h02f8: color = 2'b11;
		14'h02f9: color = 2'b11;
		14'h02fa: color = 2'b11;
		14'h02fb: color = 2'b11;
		14'h02fc: color = 2'b11;
		14'h02fd: color = 2'b11;
		14'h02fe: color = 2'b11;
		14'h02ff: color = 2'b11;
		14'h0300: color = 2'b11;
		14'h0301: color = 2'b11;
		14'h0302: color = 2'b11;
		14'h0303: color = 2'b11;
		14'h0304: color = 2'b11;
		14'h0305: color = 2'b11;
		14'h0306: color = 2'b11;
		14'h0307: color = 2'b11;
		14'h0308: color = 2'b11;
		14'h0309: color = 2'b11;
		14'h030a: color = 2'b11;
		14'h030b: color = 2'b11;
		14'h030c: color = 2'b11;
		14'h030d: color = 2'b11;
		14'h030e: color = 2'b11;
		14'h030f: color = 2'b11;
		14'h0310: color = 2'b11;
		14'h0311: color = 2'b11;
		14'h0312: color = 2'b11;
		14'h0313: color = 2'b11;
		14'h0314: color = 2'b11;
		14'h0315: color = 2'b11;
		14'h0316: color = 2'b11;
		14'h0317: color = 2'b11;
		14'h0318: color = 2'b11;
		14'h0319: color = 2'b11;
		14'h031a: color = 2'b11;
		14'h031b: color = 2'b11;
		14'h031c: color = 2'b11;
		14'h031d: color = 2'b11;
		14'h031e: color = 2'b11;
		14'h031f: color = 2'b11;
		14'h0320: color = 2'b11;
		14'h0321: color = 2'b11;
		14'h0322: color = 2'b11;
		14'h0323: color = 2'b11;
		14'h0324: color = 2'b11;
		14'h0325: color = 2'b11;
		14'h0326: color = 2'b11;
		14'h0327: color = 2'b11;
		14'h0328: color = 2'b11;
		14'h0329: color = 2'b11;
		14'h032a: color = 2'b11;
		14'h032b: color = 2'b11;
		14'h032c: color = 2'b11;
		14'h032d: color = 2'b11;
		14'h032e: color = 2'b11;
		14'h032f: color = 2'b11;
		14'h0330: color = 2'b11;
		14'h0331: color = 2'b11;
		14'h0332: color = 2'b11;
		14'h0333: color = 2'b11;
		14'h0334: color = 2'b11;
		14'h0335: color = 2'b11;
		14'h0336: color = 2'b11;
		14'h0337: color = 2'b11;
		14'h0338: color = 2'b11;
		14'h0339: color = 2'b11;
		14'h033a: color = 2'b11;
		14'h033b: color = 2'b11;
		14'h033c: color = 2'b10;
		14'h033d: color = 2'b11;
		14'h033e: color = 2'b11;
		14'h033f: color = 2'b10;
		14'h0340: color = 2'b01;
		14'h0341: color = 2'b00;
		14'h0342: color = 2'b00;
		14'h0343: color = 2'b00;
		14'h0344: color = 2'b00;
		14'h0345: color = 2'b00;
		14'h0346: color = 2'b00;
		14'h0347: color = 2'b00;
		14'h0348: color = 2'b00;
		14'h0349: color = 2'b00;
		14'h034a: color = 2'b00;
		14'h034b: color = 2'b00;
		14'h034c: color = 2'b01;
		14'h034d: color = 2'b00;
		14'h034e: color = 2'b00;
		14'h034f: color = 2'b00;
		14'h0350: color = 2'b10;
		14'h0351: color = 2'b01;
		14'h0352: color = 2'b11;
		14'h0353: color = 2'b11;
		14'h0354: color = 2'b11;
		14'h0355: color = 2'b11;
		14'h0356: color = 2'b11;
		14'h0357: color = 2'b11;
		14'h0358: color = 2'b11;
		14'h0359: color = 2'b11;
		14'h035a: color = 2'b11;
		14'h035b: color = 2'b11;
		14'h035c: color = 2'b11;
		14'h035d: color = 2'b11;
		14'h035e: color = 2'b11;
		14'h035f: color = 2'b11;
		14'h0360: color = 2'b11;
		14'h0361: color = 2'b11;
		14'h0362: color = 2'b11;
		14'h0363: color = 2'b11;
		14'h0364: color = 2'b11;
		14'h0365: color = 2'b11;
		14'h0366: color = 2'b11;
		14'h0367: color = 2'b11;
		14'h0368: color = 2'b11;
		14'h0369: color = 2'b11;
		14'h036a: color = 2'b11;
		14'h036b: color = 2'b11;
		14'h036c: color = 2'b11;
		14'h036d: color = 2'b11;
		14'h036e: color = 2'b11;
		14'h036f: color = 2'b11;
		14'h0370: color = 2'b11;
		14'h0371: color = 2'b11;
		14'h0372: color = 2'b11;
		14'h0373: color = 2'b11;
		14'h0374: color = 2'b11;
		14'h0375: color = 2'b11;
		14'h0376: color = 2'b11;
		14'h0377: color = 2'b11;
		14'h0378: color = 2'b11;
		14'h0379: color = 2'b11;
		14'h037a: color = 2'b11;
		14'h037b: color = 2'b11;
		14'h037c: color = 2'b11;
		14'h037d: color = 2'b11;
		14'h037e: color = 2'b11;
		14'h037f: color = 2'b11;
		14'h0380: color = 2'b11;
		14'h0381: color = 2'b11;
		14'h0382: color = 2'b11;
		14'h0383: color = 2'b11;
		14'h0384: color = 2'b11;
		14'h0385: color = 2'b11;
		14'h0386: color = 2'b11;
		14'h0387: color = 2'b11;
		14'h0388: color = 2'b11;
		14'h0389: color = 2'b11;
		14'h038a: color = 2'b11;
		14'h038b: color = 2'b11;
		14'h038c: color = 2'b11;
		14'h038d: color = 2'b11;
		14'h038e: color = 2'b11;
		14'h038f: color = 2'b11;
		14'h0390: color = 2'b11;
		14'h0391: color = 2'b11;
		14'h0392: color = 2'b11;
		14'h0393: color = 2'b11;
		14'h0394: color = 2'b11;
		14'h0395: color = 2'b11;
		14'h0396: color = 2'b11;
		14'h0397: color = 2'b11;
		14'h0398: color = 2'b11;
		14'h0399: color = 2'b11;
		14'h039a: color = 2'b11;
		14'h039b: color = 2'b11;
		14'h039c: color = 2'b11;
		14'h039d: color = 2'b11;
		14'h039e: color = 2'b11;
		14'h039f: color = 2'b11;
		14'h03a0: color = 2'b11;
		14'h03a1: color = 2'b11;
		14'h03a2: color = 2'b11;
		14'h03a3: color = 2'b11;
		14'h03a4: color = 2'b11;
		14'h03a5: color = 2'b11;
		14'h03a6: color = 2'b11;
		14'h03a7: color = 2'b11;
		14'h03a8: color = 2'b11;
		14'h03a9: color = 2'b11;
		14'h03aa: color = 2'b11;
		14'h03ab: color = 2'b11;
		14'h03ac: color = 2'b11;
		14'h03ad: color = 2'b11;
		14'h03ae: color = 2'b11;
		14'h03af: color = 2'b11;
		14'h03b0: color = 2'b11;
		14'h03b1: color = 2'b11;
		14'h03b2: color = 2'b11;
		14'h03b3: color = 2'b11;
		14'h03b4: color = 2'b11;
		14'h03b5: color = 2'b11;
		14'h03b6: color = 2'b11;
		14'h03b7: color = 2'b11;
		14'h03b8: color = 2'b11;
		14'h03b9: color = 2'b10;
		14'h03ba: color = 2'b10;
		14'h03bb: color = 2'b01;
		14'h03bc: color = 2'b00;
		14'h03bd: color = 2'b00;
		14'h03be: color = 2'b01;
		14'h03bf: color = 2'b01;
		14'h03c0: color = 2'b00;
		14'h03c1: color = 2'b00;
		14'h03c2: color = 2'b00;
		14'h03c3: color = 2'b00;
		14'h03c4: color = 2'b00;
		14'h03c5: color = 2'b00;
		14'h03c6: color = 2'b00;
		14'h03c7: color = 2'b00;
		14'h03c8: color = 2'b00;
		14'h03c9: color = 2'b00;
		14'h03ca: color = 2'b00;
		14'h03cb: color = 2'b00;
		14'h03cc: color = 2'b00;
		14'h03cd: color = 2'b00;
		14'h03ce: color = 2'b00;
		14'h03cf: color = 2'b00;
		14'h03d0: color = 2'b00;
		14'h03d1: color = 2'b00;
		14'h03d2: color = 2'b00;
		14'h03d3: color = 2'b01;
		14'h03d4: color = 2'b01;
		14'h03d5: color = 2'b11;
		14'h03d6: color = 2'b11;
		14'h03d7: color = 2'b11;
		14'h03d8: color = 2'b11;
		14'h03d9: color = 2'b11;
		14'h03da: color = 2'b11;
		14'h03db: color = 2'b11;
		14'h03dc: color = 2'b11;
		14'h03dd: color = 2'b11;
		14'h03de: color = 2'b11;
		14'h03df: color = 2'b11;
		14'h03e0: color = 2'b11;
		14'h03e1: color = 2'b11;
		14'h03e2: color = 2'b11;
		14'h03e3: color = 2'b11;
		14'h03e4: color = 2'b11;
		14'h03e5: color = 2'b11;
		14'h03e6: color = 2'b11;
		14'h03e7: color = 2'b11;
		14'h03e8: color = 2'b11;
		14'h03e9: color = 2'b11;
		14'h03ea: color = 2'b11;
		14'h03eb: color = 2'b11;
		14'h03ec: color = 2'b11;
		14'h03ed: color = 2'b11;
		14'h03ee: color = 2'b11;
		14'h03ef: color = 2'b11;
		14'h03f0: color = 2'b11;
		14'h03f1: color = 2'b11;
		14'h03f2: color = 2'b11;
		14'h03f3: color = 2'b11;
		14'h03f4: color = 2'b11;
		14'h03f5: color = 2'b11;
		14'h03f6: color = 2'b11;
		14'h03f7: color = 2'b11;
		14'h03f8: color = 2'b11;
		14'h03f9: color = 2'b11;
		14'h03fa: color = 2'b11;
		14'h03fb: color = 2'b11;
		14'h03fc: color = 2'b11;
		14'h03fd: color = 2'b11;
		14'h03fe: color = 2'b11;
		14'h03ff: color = 2'b11;
		14'h0400: color = 2'b11;
		14'h0401: color = 2'b11;
		14'h0402: color = 2'b11;
		14'h0403: color = 2'b11;
		14'h0404: color = 2'b11;
		14'h0405: color = 2'b11;
		14'h0406: color = 2'b11;
		14'h0407: color = 2'b11;
		14'h0408: color = 2'b11;
		14'h0409: color = 2'b11;
		14'h040a: color = 2'b11;
		14'h040b: color = 2'b11;
		14'h040c: color = 2'b11;
		14'h040d: color = 2'b11;
		14'h040e: color = 2'b11;
		14'h040f: color = 2'b11;
		14'h0410: color = 2'b11;
		14'h0411: color = 2'b11;
		14'h0412: color = 2'b11;
		14'h0413: color = 2'b11;
		14'h0414: color = 2'b11;
		14'h0415: color = 2'b11;
		14'h0416: color = 2'b11;
		14'h0417: color = 2'b11;
		14'h0418: color = 2'b11;
		14'h0419: color = 2'b11;
		14'h041a: color = 2'b11;
		14'h041b: color = 2'b11;
		14'h041c: color = 2'b11;
		14'h041d: color = 2'b11;
		14'h041e: color = 2'b11;
		14'h041f: color = 2'b11;
		14'h0420: color = 2'b11;
		14'h0421: color = 2'b11;
		14'h0422: color = 2'b11;
		14'h0423: color = 2'b11;
		14'h0424: color = 2'b11;
		14'h0425: color = 2'b11;
		14'h0426: color = 2'b11;
		14'h0427: color = 2'b11;
		14'h0428: color = 2'b11;
		14'h0429: color = 2'b11;
		14'h042a: color = 2'b11;
		14'h042b: color = 2'b11;
		14'h042c: color = 2'b11;
		14'h042d: color = 2'b11;
		14'h042e: color = 2'b11;
		14'h042f: color = 2'b11;
		14'h0430: color = 2'b11;
		14'h0431: color = 2'b11;
		14'h0432: color = 2'b11;
		14'h0433: color = 2'b11;
		14'h0434: color = 2'b11;
		14'h0435: color = 2'b11;
		14'h0436: color = 2'b11;
		14'h0437: color = 2'b11;
		14'h0438: color = 2'b11;
		14'h0439: color = 2'b10;
		14'h043a: color = 2'b10;
		14'h043b: color = 2'b01;
		14'h043c: color = 2'b00;
		14'h043d: color = 2'b00;
		14'h043e: color = 2'b01;
		14'h043f: color = 2'b01;
		14'h0440: color = 2'b00;
		14'h0441: color = 2'b00;
		14'h0442: color = 2'b00;
		14'h0443: color = 2'b00;
		14'h0444: color = 2'b00;
		14'h0445: color = 2'b00;
		14'h0446: color = 2'b00;
		14'h0447: color = 2'b00;
		14'h0448: color = 2'b00;
		14'h0449: color = 2'b00;
		14'h044a: color = 2'b00;
		14'h044b: color = 2'b00;
		14'h044c: color = 2'b00;
		14'h044d: color = 2'b00;
		14'h044e: color = 2'b00;
		14'h044f: color = 2'b00;
		14'h0450: color = 2'b00;
		14'h0451: color = 2'b00;
		14'h0452: color = 2'b00;
		14'h0453: color = 2'b01;
		14'h0454: color = 2'b01;
		14'h0455: color = 2'b11;
		14'h0456: color = 2'b11;
		14'h0457: color = 2'b11;
		14'h0458: color = 2'b11;
		14'h0459: color = 2'b11;
		14'h045a: color = 2'b11;
		14'h045b: color = 2'b11;
		14'h045c: color = 2'b11;
		14'h045d: color = 2'b11;
		14'h045e: color = 2'b11;
		14'h045f: color = 2'b11;
		14'h0460: color = 2'b11;
		14'h0461: color = 2'b11;
		14'h0462: color = 2'b11;
		14'h0463: color = 2'b11;
		14'h0464: color = 2'b11;
		14'h0465: color = 2'b11;
		14'h0466: color = 2'b11;
		14'h0467: color = 2'b11;
		14'h0468: color = 2'b11;
		14'h0469: color = 2'b11;
		14'h046a: color = 2'b11;
		14'h046b: color = 2'b11;
		14'h046c: color = 2'b11;
		14'h046d: color = 2'b11;
		14'h046e: color = 2'b11;
		14'h046f: color = 2'b11;
		14'h0470: color = 2'b11;
		14'h0471: color = 2'b11;
		14'h0472: color = 2'b11;
		14'h0473: color = 2'b11;
		14'h0474: color = 2'b11;
		14'h0475: color = 2'b11;
		14'h0476: color = 2'b11;
		14'h0477: color = 2'b11;
		14'h0478: color = 2'b11;
		14'h0479: color = 2'b11;
		14'h047a: color = 2'b11;
		14'h047b: color = 2'b11;
		14'h047c: color = 2'b11;
		14'h047d: color = 2'b11;
		14'h047e: color = 2'b11;
		14'h047f: color = 2'b11;
		14'h0480: color = 2'b11;
		14'h0481: color = 2'b11;
		14'h0482: color = 2'b11;
		14'h0483: color = 2'b11;
		14'h0484: color = 2'b11;
		14'h0485: color = 2'b11;
		14'h0486: color = 2'b11;
		14'h0487: color = 2'b11;
		14'h0488: color = 2'b11;
		14'h0489: color = 2'b11;
		14'h048a: color = 2'b11;
		14'h048b: color = 2'b11;
		14'h048c: color = 2'b11;
		14'h048d: color = 2'b11;
		14'h048e: color = 2'b11;
		14'h048f: color = 2'b11;
		14'h0490: color = 2'b11;
		14'h0491: color = 2'b11;
		14'h0492: color = 2'b11;
		14'h0493: color = 2'b11;
		14'h0494: color = 2'b11;
		14'h0495: color = 2'b11;
		14'h0496: color = 2'b11;
		14'h0497: color = 2'b11;
		14'h0498: color = 2'b11;
		14'h0499: color = 2'b11;
		14'h049a: color = 2'b11;
		14'h049b: color = 2'b11;
		14'h049c: color = 2'b11;
		14'h049d: color = 2'b11;
		14'h049e: color = 2'b11;
		14'h049f: color = 2'b11;
		14'h04a0: color = 2'b11;
		14'h04a1: color = 2'b11;
		14'h04a2: color = 2'b11;
		14'h04a3: color = 2'b11;
		14'h04a4: color = 2'b11;
		14'h04a5: color = 2'b11;
		14'h04a6: color = 2'b11;
		14'h04a7: color = 2'b11;
		14'h04a8: color = 2'b11;
		14'h04a9: color = 2'b11;
		14'h04aa: color = 2'b11;
		14'h04ab: color = 2'b11;
		14'h04ac: color = 2'b11;
		14'h04ad: color = 2'b11;
		14'h04ae: color = 2'b11;
		14'h04af: color = 2'b11;
		14'h04b0: color = 2'b11;
		14'h04b1: color = 2'b11;
		14'h04b2: color = 2'b11;
		14'h04b3: color = 2'b11;
		14'h04b4: color = 2'b11;
		14'h04b5: color = 2'b11;
		14'h04b6: color = 2'b10;
		14'h04b7: color = 2'b10;
		14'h04b8: color = 2'b10;
		14'h04b9: color = 2'b01;
		14'h04ba: color = 2'b00;
		14'h04bb: color = 2'b00;
		14'h04bc: color = 2'b01;
		14'h04bd: color = 2'b01;
		14'h04be: color = 2'b00;
		14'h04bf: color = 2'b01;
		14'h04c0: color = 2'b01;
		14'h04c1: color = 2'b01;
		14'h04c2: color = 2'b00;
		14'h04c3: color = 2'b01;
		14'h04c4: color = 2'b00;
		14'h04c5: color = 2'b01;
		14'h04c6: color = 2'b00;
		14'h04c7: color = 2'b00;
		14'h04c8: color = 2'b00;
		14'h04c9: color = 2'b01;
		14'h04ca: color = 2'b00;
		14'h04cb: color = 2'b00;
		14'h04cc: color = 2'b00;
		14'h04cd: color = 2'b00;
		14'h04ce: color = 2'b00;
		14'h04cf: color = 2'b00;
		14'h04d0: color = 2'b00;
		14'h04d1: color = 2'b00;
		14'h04d2: color = 2'b00;
		14'h04d3: color = 2'b00;
		14'h04d4: color = 2'b00;
		14'h04d5: color = 2'b00;
		14'h04d6: color = 2'b00;
		14'h04d7: color = 2'b11;
		14'h04d8: color = 2'b11;
		14'h04d9: color = 2'b11;
		14'h04da: color = 2'b11;
		14'h04db: color = 2'b11;
		14'h04dc: color = 2'b11;
		14'h04dd: color = 2'b11;
		14'h04de: color = 2'b11;
		14'h04df: color = 2'b11;
		14'h04e0: color = 2'b11;
		14'h04e1: color = 2'b11;
		14'h04e2: color = 2'b11;
		14'h04e3: color = 2'b11;
		14'h04e4: color = 2'b11;
		14'h04e5: color = 2'b11;
		14'h04e6: color = 2'b11;
		14'h04e7: color = 2'b11;
		14'h04e8: color = 2'b11;
		14'h04e9: color = 2'b11;
		14'h04ea: color = 2'b11;
		14'h04eb: color = 2'b11;
		14'h04ec: color = 2'b11;
		14'h04ed: color = 2'b11;
		14'h04ee: color = 2'b11;
		14'h04ef: color = 2'b11;
		14'h04f0: color = 2'b11;
		14'h04f1: color = 2'b11;
		14'h04f2: color = 2'b11;
		14'h04f3: color = 2'b11;
		14'h04f4: color = 2'b11;
		14'h04f5: color = 2'b11;
		14'h04f6: color = 2'b11;
		14'h04f7: color = 2'b11;
		14'h04f8: color = 2'b11;
		14'h04f9: color = 2'b11;
		14'h04fa: color = 2'b11;
		14'h04fb: color = 2'b11;
		14'h04fc: color = 2'b11;
		14'h04fd: color = 2'b11;
		14'h04fe: color = 2'b11;
		14'h04ff: color = 2'b11;
		14'h0500: color = 2'b11;
		14'h0501: color = 2'b11;
		14'h0502: color = 2'b11;
		14'h0503: color = 2'b11;
		14'h0504: color = 2'b11;
		14'h0505: color = 2'b11;
		14'h0506: color = 2'b11;
		14'h0507: color = 2'b11;
		14'h0508: color = 2'b11;
		14'h0509: color = 2'b11;
		14'h050a: color = 2'b11;
		14'h050b: color = 2'b11;
		14'h050c: color = 2'b11;
		14'h050d: color = 2'b11;
		14'h050e: color = 2'b11;
		14'h050f: color = 2'b11;
		14'h0510: color = 2'b11;
		14'h0511: color = 2'b11;
		14'h0512: color = 2'b11;
		14'h0513: color = 2'b11;
		14'h0514: color = 2'b11;
		14'h0515: color = 2'b11;
		14'h0516: color = 2'b11;
		14'h0517: color = 2'b11;
		14'h0518: color = 2'b11;
		14'h0519: color = 2'b11;
		14'h051a: color = 2'b11;
		14'h051b: color = 2'b11;
		14'h051c: color = 2'b11;
		14'h051d: color = 2'b11;
		14'h051e: color = 2'b11;
		14'h051f: color = 2'b11;
		14'h0520: color = 2'b11;
		14'h0521: color = 2'b11;
		14'h0522: color = 2'b11;
		14'h0523: color = 2'b11;
		14'h0524: color = 2'b11;
		14'h0525: color = 2'b11;
		14'h0526: color = 2'b11;
		14'h0527: color = 2'b11;
		14'h0528: color = 2'b11;
		14'h0529: color = 2'b11;
		14'h052a: color = 2'b11;
		14'h052b: color = 2'b11;
		14'h052c: color = 2'b11;
		14'h052d: color = 2'b11;
		14'h052e: color = 2'b11;
		14'h052f: color = 2'b11;
		14'h0530: color = 2'b11;
		14'h0531: color = 2'b11;
		14'h0532: color = 2'b11;
		14'h0533: color = 2'b10;
		14'h0534: color = 2'b01;
		14'h0535: color = 2'b00;
		14'h0536: color = 2'b01;
		14'h0537: color = 2'b01;
		14'h0538: color = 2'b01;
		14'h0539: color = 2'b01;
		14'h053a: color = 2'b01;
		14'h053b: color = 2'b01;
		14'h053c: color = 2'b00;
		14'h053d: color = 2'b01;
		14'h053e: color = 2'b01;
		14'h053f: color = 2'b00;
		14'h0540: color = 2'b00;
		14'h0541: color = 2'b00;
		14'h0542: color = 2'b01;
		14'h0543: color = 2'b00;
		14'h0544: color = 2'b00;
		14'h0545: color = 2'b01;
		14'h0546: color = 2'b01;
		14'h0547: color = 2'b00;
		14'h0548: color = 2'b00;
		14'h0549: color = 2'b00;
		14'h054a: color = 2'b00;
		14'h054b: color = 2'b00;
		14'h054c: color = 2'b00;
		14'h054d: color = 2'b00;
		14'h054e: color = 2'b00;
		14'h054f: color = 2'b00;
		14'h0550: color = 2'b00;
		14'h0551: color = 2'b00;
		14'h0552: color = 2'b00;
		14'h0553: color = 2'b00;
		14'h0554: color = 2'b00;
		14'h0555: color = 2'b00;
		14'h0556: color = 2'b00;
		14'h0557: color = 2'b00;
		14'h0558: color = 2'b00;
		14'h0559: color = 2'b00;
		14'h055a: color = 2'b11;
		14'h055b: color = 2'b11;
		14'h055c: color = 2'b11;
		14'h055d: color = 2'b11;
		14'h055e: color = 2'b11;
		14'h055f: color = 2'b11;
		14'h0560: color = 2'b11;
		14'h0561: color = 2'b11;
		14'h0562: color = 2'b11;
		14'h0563: color = 2'b11;
		14'h0564: color = 2'b11;
		14'h0565: color = 2'b11;
		14'h0566: color = 2'b11;
		14'h0567: color = 2'b11;
		14'h0568: color = 2'b11;
		14'h0569: color = 2'b11;
		14'h056a: color = 2'b11;
		14'h056b: color = 2'b11;
		14'h056c: color = 2'b11;
		14'h056d: color = 2'b11;
		14'h056e: color = 2'b11;
		14'h056f: color = 2'b11;
		14'h0570: color = 2'b11;
		14'h0571: color = 2'b11;
		14'h0572: color = 2'b11;
		14'h0573: color = 2'b11;
		14'h0574: color = 2'b11;
		14'h0575: color = 2'b11;
		14'h0576: color = 2'b11;
		14'h0577: color = 2'b11;
		14'h0578: color = 2'b11;
		14'h0579: color = 2'b11;
		14'h057a: color = 2'b11;
		14'h057b: color = 2'b11;
		14'h057c: color = 2'b11;
		14'h057d: color = 2'b11;
		14'h057e: color = 2'b11;
		14'h057f: color = 2'b11;
		14'h0580: color = 2'b11;
		14'h0581: color = 2'b11;
		14'h0582: color = 2'b11;
		14'h0583: color = 2'b11;
		14'h0584: color = 2'b11;
		14'h0585: color = 2'b11;
		14'h0586: color = 2'b11;
		14'h0587: color = 2'b11;
		14'h0588: color = 2'b11;
		14'h0589: color = 2'b11;
		14'h058a: color = 2'b11;
		14'h058b: color = 2'b11;
		14'h058c: color = 2'b11;
		14'h058d: color = 2'b11;
		14'h058e: color = 2'b11;
		14'h058f: color = 2'b11;
		14'h0590: color = 2'b11;
		14'h0591: color = 2'b11;
		14'h0592: color = 2'b11;
		14'h0593: color = 2'b11;
		14'h0594: color = 2'b11;
		14'h0595: color = 2'b11;
		14'h0596: color = 2'b11;
		14'h0597: color = 2'b11;
		14'h0598: color = 2'b11;
		14'h0599: color = 2'b11;
		14'h059a: color = 2'b11;
		14'h059b: color = 2'b11;
		14'h059c: color = 2'b11;
		14'h059d: color = 2'b11;
		14'h059e: color = 2'b11;
		14'h059f: color = 2'b11;
		14'h05a0: color = 2'b11;
		14'h05a1: color = 2'b11;
		14'h05a2: color = 2'b11;
		14'h05a3: color = 2'b11;
		14'h05a4: color = 2'b11;
		14'h05a5: color = 2'b11;
		14'h05a6: color = 2'b11;
		14'h05a7: color = 2'b11;
		14'h05a8: color = 2'b11;
		14'h05a9: color = 2'b11;
		14'h05aa: color = 2'b11;
		14'h05ab: color = 2'b11;
		14'h05ac: color = 2'b11;
		14'h05ad: color = 2'b11;
		14'h05ae: color = 2'b11;
		14'h05af: color = 2'b11;
		14'h05b0: color = 2'b11;
		14'h05b1: color = 2'b11;
		14'h05b2: color = 2'b10;
		14'h05b3: color = 2'b11;
		14'h05b4: color = 2'b01;
		14'h05b5: color = 2'b00;
		14'h05b6: color = 2'b01;
		14'h05b7: color = 2'b00;
		14'h05b8: color = 2'b00;
		14'h05b9: color = 2'b00;
		14'h05ba: color = 2'b00;
		14'h05bb: color = 2'b00;
		14'h05bc: color = 2'b00;
		14'h05bd: color = 2'b01;
		14'h05be: color = 2'b01;
		14'h05bf: color = 2'b01;
		14'h05c0: color = 2'b01;
		14'h05c1: color = 2'b01;
		14'h05c2: color = 2'b01;
		14'h05c3: color = 2'b01;
		14'h05c4: color = 2'b00;
		14'h05c5: color = 2'b01;
		14'h05c6: color = 2'b00;
		14'h05c7: color = 2'b01;
		14'h05c8: color = 2'b01;
		14'h05c9: color = 2'b00;
		14'h05ca: color = 2'b00;
		14'h05cb: color = 2'b00;
		14'h05cc: color = 2'b00;
		14'h05cd: color = 2'b00;
		14'h05ce: color = 2'b00;
		14'h05cf: color = 2'b00;
		14'h05d0: color = 2'b00;
		14'h05d1: color = 2'b00;
		14'h05d2: color = 2'b00;
		14'h05d3: color = 2'b00;
		14'h05d4: color = 2'b00;
		14'h05d5: color = 2'b00;
		14'h05d6: color = 2'b00;
		14'h05d7: color = 2'b00;
		14'h05d8: color = 2'b00;
		14'h05d9: color = 2'b00;
		14'h05da: color = 2'b00;
		14'h05db: color = 2'b01;
		14'h05dc: color = 2'b10;
		14'h05dd: color = 2'b11;
		14'h05de: color = 2'b11;
		14'h05df: color = 2'b11;
		14'h05e0: color = 2'b11;
		14'h05e1: color = 2'b11;
		14'h05e2: color = 2'b11;
		14'h05e3: color = 2'b11;
		14'h05e4: color = 2'b11;
		14'h05e5: color = 2'b11;
		14'h05e6: color = 2'b11;
		14'h05e7: color = 2'b11;
		14'h05e8: color = 2'b11;
		14'h05e9: color = 2'b11;
		14'h05ea: color = 2'b11;
		14'h05eb: color = 2'b11;
		14'h05ec: color = 2'b11;
		14'h05ed: color = 2'b11;
		14'h05ee: color = 2'b11;
		14'h05ef: color = 2'b11;
		14'h05f0: color = 2'b11;
		14'h05f1: color = 2'b11;
		14'h05f2: color = 2'b11;
		14'h05f3: color = 2'b11;
		14'h05f4: color = 2'b11;
		14'h05f5: color = 2'b11;
		14'h05f6: color = 2'b11;
		14'h05f7: color = 2'b11;
		14'h05f8: color = 2'b11;
		14'h05f9: color = 2'b11;
		14'h05fa: color = 2'b11;
		14'h05fb: color = 2'b11;
		14'h05fc: color = 2'b11;
		14'h05fd: color = 2'b11;
		14'h05fe: color = 2'b11;
		14'h05ff: color = 2'b11;
		14'h0600: color = 2'b11;
		14'h0601: color = 2'b11;
		14'h0602: color = 2'b11;
		14'h0603: color = 2'b11;
		14'h0604: color = 2'b11;
		14'h0605: color = 2'b11;
		14'h0606: color = 2'b11;
		14'h0607: color = 2'b11;
		14'h0608: color = 2'b11;
		14'h0609: color = 2'b11;
		14'h060a: color = 2'b11;
		14'h060b: color = 2'b11;
		14'h060c: color = 2'b11;
		14'h060d: color = 2'b11;
		14'h060e: color = 2'b11;
		14'h060f: color = 2'b11;
		14'h0610: color = 2'b11;
		14'h0611: color = 2'b11;
		14'h0612: color = 2'b11;
		14'h0613: color = 2'b11;
		14'h0614: color = 2'b11;
		14'h0615: color = 2'b11;
		14'h0616: color = 2'b11;
		14'h0617: color = 2'b11;
		14'h0618: color = 2'b11;
		14'h0619: color = 2'b11;
		14'h061a: color = 2'b11;
		14'h061b: color = 2'b11;
		14'h061c: color = 2'b11;
		14'h061d: color = 2'b11;
		14'h061e: color = 2'b11;
		14'h061f: color = 2'b11;
		14'h0620: color = 2'b11;
		14'h0621: color = 2'b11;
		14'h0622: color = 2'b11;
		14'h0623: color = 2'b11;
		14'h0624: color = 2'b11;
		14'h0625: color = 2'b11;
		14'h0626: color = 2'b11;
		14'h0627: color = 2'b11;
		14'h0628: color = 2'b11;
		14'h0629: color = 2'b11;
		14'h062a: color = 2'b11;
		14'h062b: color = 2'b11;
		14'h062c: color = 2'b11;
		14'h062d: color = 2'b11;
		14'h062e: color = 2'b11;
		14'h062f: color = 2'b11;
		14'h0630: color = 2'b11;
		14'h0631: color = 2'b11;
		14'h0632: color = 2'b10;
		14'h0633: color = 2'b01;
		14'h0634: color = 2'b00;
		14'h0635: color = 2'b00;
		14'h0636: color = 2'b00;
		14'h0637: color = 2'b00;
		14'h0638: color = 2'b00;
		14'h0639: color = 2'b00;
		14'h063a: color = 2'b00;
		14'h063b: color = 2'b00;
		14'h063c: color = 2'b00;
		14'h063d: color = 2'b01;
		14'h063e: color = 2'b01;
		14'h063f: color = 2'b01;
		14'h0640: color = 2'b00;
		14'h0641: color = 2'b01;
		14'h0642: color = 2'b00;
		14'h0643: color = 2'b00;
		14'h0644: color = 2'b00;
		14'h0645: color = 2'b00;
		14'h0646: color = 2'b00;
		14'h0647: color = 2'b01;
		14'h0648: color = 2'b01;
		14'h0649: color = 2'b00;
		14'h064a: color = 2'b01;
		14'h064b: color = 2'b00;
		14'h064c: color = 2'b00;
		14'h064d: color = 2'b00;
		14'h064e: color = 2'b00;
		14'h064f: color = 2'b00;
		14'h0650: color = 2'b00;
		14'h0651: color = 2'b00;
		14'h0652: color = 2'b00;
		14'h0653: color = 2'b00;
		14'h0654: color = 2'b00;
		14'h0655: color = 2'b00;
		14'h0656: color = 2'b00;
		14'h0657: color = 2'b00;
		14'h0658: color = 2'b00;
		14'h0659: color = 2'b00;
		14'h065a: color = 2'b00;
		14'h065b: color = 2'b00;
		14'h065c: color = 2'b00;
		14'h065d: color = 2'b01;
		14'h065e: color = 2'b11;
		14'h065f: color = 2'b11;
		14'h0660: color = 2'b11;
		14'h0661: color = 2'b11;
		14'h0662: color = 2'b11;
		14'h0663: color = 2'b11;
		14'h0664: color = 2'b11;
		14'h0665: color = 2'b11;
		14'h0666: color = 2'b11;
		14'h0667: color = 2'b11;
		14'h0668: color = 2'b11;
		14'h0669: color = 2'b11;
		14'h066a: color = 2'b11;
		14'h066b: color = 2'b11;
		14'h066c: color = 2'b11;
		14'h066d: color = 2'b11;
		14'h066e: color = 2'b11;
		14'h066f: color = 2'b11;
		14'h0670: color = 2'b11;
		14'h0671: color = 2'b11;
		14'h0672: color = 2'b11;
		14'h0673: color = 2'b11;
		14'h0674: color = 2'b11;
		14'h0675: color = 2'b11;
		14'h0676: color = 2'b11;
		14'h0677: color = 2'b11;
		14'h0678: color = 2'b11;
		14'h0679: color = 2'b11;
		14'h067a: color = 2'b11;
		14'h067b: color = 2'b11;
		14'h067c: color = 2'b11;
		14'h067d: color = 2'b11;
		14'h067e: color = 2'b11;
		14'h067f: color = 2'b11;
		14'h0680: color = 2'b11;
		14'h0681: color = 2'b11;
		14'h0682: color = 2'b11;
		14'h0683: color = 2'b11;
		14'h0684: color = 2'b11;
		14'h0685: color = 2'b11;
		14'h0686: color = 2'b11;
		14'h0687: color = 2'b11;
		14'h0688: color = 2'b11;
		14'h0689: color = 2'b11;
		14'h068a: color = 2'b11;
		14'h068b: color = 2'b11;
		14'h068c: color = 2'b11;
		14'h068d: color = 2'b11;
		14'h068e: color = 2'b11;
		14'h068f: color = 2'b11;
		14'h0690: color = 2'b11;
		14'h0691: color = 2'b11;
		14'h0692: color = 2'b11;
		14'h0693: color = 2'b11;
		14'h0694: color = 2'b11;
		14'h0695: color = 2'b11;
		14'h0696: color = 2'b11;
		14'h0697: color = 2'b11;
		14'h0698: color = 2'b11;
		14'h0699: color = 2'b11;
		14'h069a: color = 2'b11;
		14'h069b: color = 2'b11;
		14'h069c: color = 2'b11;
		14'h069d: color = 2'b11;
		14'h069e: color = 2'b11;
		14'h069f: color = 2'b11;
		14'h06a0: color = 2'b11;
		14'h06a1: color = 2'b11;
		14'h06a2: color = 2'b11;
		14'h06a3: color = 2'b11;
		14'h06a4: color = 2'b11;
		14'h06a5: color = 2'b11;
		14'h06a6: color = 2'b11;
		14'h06a7: color = 2'b11;
		14'h06a8: color = 2'b11;
		14'h06a9: color = 2'b11;
		14'h06aa: color = 2'b11;
		14'h06ab: color = 2'b11;
		14'h06ac: color = 2'b11;
		14'h06ad: color = 2'b11;
		14'h06ae: color = 2'b01;
		14'h06af: color = 2'b00;
		14'h06b0: color = 2'b01;
		14'h06b1: color = 2'b11;
		14'h06b2: color = 2'b01;
		14'h06b3: color = 2'b00;
		14'h06b4: color = 2'b00;
		14'h06b5: color = 2'b00;
		14'h06b6: color = 2'b00;
		14'h06b7: color = 2'b00;
		14'h06b8: color = 2'b00;
		14'h06b9: color = 2'b00;
		14'h06ba: color = 2'b00;
		14'h06bb: color = 2'b01;
		14'h06bc: color = 2'b01;
		14'h06bd: color = 2'b00;
		14'h06be: color = 2'b00;
		14'h06bf: color = 2'b00;
		14'h06c0: color = 2'b00;
		14'h06c1: color = 2'b00;
		14'h06c2: color = 2'b01;
		14'h06c3: color = 2'b00;
		14'h06c4: color = 2'b00;
		14'h06c5: color = 2'b00;
		14'h06c6: color = 2'b01;
		14'h06c7: color = 2'b00;
		14'h06c8: color = 2'b00;
		14'h06c9: color = 2'b01;
		14'h06ca: color = 2'b01;
		14'h06cb: color = 2'b00;
		14'h06cc: color = 2'b00;
		14'h06cd: color = 2'b00;
		14'h06ce: color = 2'b00;
		14'h06cf: color = 2'b00;
		14'h06d0: color = 2'b00;
		14'h06d1: color = 2'b00;
		14'h06d2: color = 2'b00;
		14'h06d3: color = 2'b00;
		14'h06d4: color = 2'b00;
		14'h06d5: color = 2'b00;
		14'h06d6: color = 2'b00;
		14'h06d7: color = 2'b00;
		14'h06d8: color = 2'b00;
		14'h06d9: color = 2'b00;
		14'h06da: color = 2'b00;
		14'h06db: color = 2'b00;
		14'h06dc: color = 2'b00;
		14'h06dd: color = 2'b00;
		14'h06de: color = 2'b00;
		14'h06df: color = 2'b10;
		14'h06e0: color = 2'b11;
		14'h06e1: color = 2'b11;
		14'h06e2: color = 2'b11;
		14'h06e3: color = 2'b11;
		14'h06e4: color = 2'b11;
		14'h06e5: color = 2'b11;
		14'h06e6: color = 2'b11;
		14'h06e7: color = 2'b11;
		14'h06e8: color = 2'b11;
		14'h06e9: color = 2'b11;
		14'h06ea: color = 2'b11;
		14'h06eb: color = 2'b11;
		14'h06ec: color = 2'b11;
		14'h06ed: color = 2'b11;
		14'h06ee: color = 2'b11;
		14'h06ef: color = 2'b11;
		14'h06f0: color = 2'b11;
		14'h06f1: color = 2'b11;
		14'h06f2: color = 2'b11;
		14'h06f3: color = 2'b11;
		14'h06f4: color = 2'b11;
		14'h06f5: color = 2'b11;
		14'h06f6: color = 2'b11;
		14'h06f7: color = 2'b11;
		14'h06f8: color = 2'b11;
		14'h06f9: color = 2'b11;
		14'h06fa: color = 2'b11;
		14'h06fb: color = 2'b11;
		14'h06fc: color = 2'b11;
		14'h06fd: color = 2'b11;
		14'h06fe: color = 2'b11;
		14'h06ff: color = 2'b11;
		14'h0700: color = 2'b11;
		14'h0701: color = 2'b11;
		14'h0702: color = 2'b11;
		14'h0703: color = 2'b11;
		14'h0704: color = 2'b11;
		14'h0705: color = 2'b11;
		14'h0706: color = 2'b11;
		14'h0707: color = 2'b11;
		14'h0708: color = 2'b11;
		14'h0709: color = 2'b11;
		14'h070a: color = 2'b11;
		14'h070b: color = 2'b11;
		14'h070c: color = 2'b11;
		14'h070d: color = 2'b11;
		14'h070e: color = 2'b11;
		14'h070f: color = 2'b11;
		14'h0710: color = 2'b11;
		14'h0711: color = 2'b11;
		14'h0712: color = 2'b11;
		14'h0713: color = 2'b11;
		14'h0714: color = 2'b11;
		14'h0715: color = 2'b11;
		14'h0716: color = 2'b11;
		14'h0717: color = 2'b11;
		14'h0718: color = 2'b11;
		14'h0719: color = 2'b11;
		14'h071a: color = 2'b11;
		14'h071b: color = 2'b11;
		14'h071c: color = 2'b11;
		14'h071d: color = 2'b11;
		14'h071e: color = 2'b11;
		14'h071f: color = 2'b11;
		14'h0720: color = 2'b11;
		14'h0721: color = 2'b11;
		14'h0722: color = 2'b11;
		14'h0723: color = 2'b11;
		14'h0724: color = 2'b11;
		14'h0725: color = 2'b11;
		14'h0726: color = 2'b11;
		14'h0727: color = 2'b11;
		14'h0728: color = 2'b11;
		14'h0729: color = 2'b11;
		14'h072a: color = 2'b11;
		14'h072b: color = 2'b11;
		14'h072c: color = 2'b10;
		14'h072d: color = 2'b00;
		14'h072e: color = 2'b00;
		14'h072f: color = 2'b00;
		14'h0730: color = 2'b01;
		14'h0731: color = 2'b01;
		14'h0732: color = 2'b00;
		14'h0733: color = 2'b00;
		14'h0734: color = 2'b00;
		14'h0735: color = 2'b00;
		14'h0736: color = 2'b00;
		14'h0737: color = 2'b00;
		14'h0738: color = 2'b00;
		14'h0739: color = 2'b00;
		14'h073a: color = 2'b00;
		14'h073b: color = 2'b00;
		14'h073c: color = 2'b01;
		14'h073d: color = 2'b00;
		14'h073e: color = 2'b00;
		14'h073f: color = 2'b00;
		14'h0740: color = 2'b00;
		14'h0741: color = 2'b00;
		14'h0742: color = 2'b00;
		14'h0743: color = 2'b00;
		14'h0744: color = 2'b00;
		14'h0745: color = 2'b00;
		14'h0746: color = 2'b00;
		14'h0747: color = 2'b00;
		14'h0748: color = 2'b00;
		14'h0749: color = 2'b00;
		14'h074a: color = 2'b00;
		14'h074b: color = 2'b00;
		14'h074c: color = 2'b00;
		14'h074d: color = 2'b00;
		14'h074e: color = 2'b00;
		14'h074f: color = 2'b00;
		14'h0750: color = 2'b00;
		14'h0751: color = 2'b00;
		14'h0752: color = 2'b00;
		14'h0753: color = 2'b00;
		14'h0754: color = 2'b00;
		14'h0755: color = 2'b00;
		14'h0756: color = 2'b00;
		14'h0757: color = 2'b00;
		14'h0758: color = 2'b00;
		14'h0759: color = 2'b00;
		14'h075a: color = 2'b00;
		14'h075b: color = 2'b00;
		14'h075c: color = 2'b00;
		14'h075d: color = 2'b00;
		14'h075e: color = 2'b00;
		14'h075f: color = 2'b00;
		14'h0760: color = 2'b10;
		14'h0761: color = 2'b11;
		14'h0762: color = 2'b11;
		14'h0763: color = 2'b11;
		14'h0764: color = 2'b11;
		14'h0765: color = 2'b11;
		14'h0766: color = 2'b11;
		14'h0767: color = 2'b11;
		14'h0768: color = 2'b11;
		14'h0769: color = 2'b11;
		14'h076a: color = 2'b11;
		14'h076b: color = 2'b11;
		14'h076c: color = 2'b11;
		14'h076d: color = 2'b11;
		14'h076e: color = 2'b11;
		14'h076f: color = 2'b11;
		14'h0770: color = 2'b11;
		14'h0771: color = 2'b11;
		14'h0772: color = 2'b11;
		14'h0773: color = 2'b11;
		14'h0774: color = 2'b11;
		14'h0775: color = 2'b11;
		14'h0776: color = 2'b11;
		14'h0777: color = 2'b11;
		14'h0778: color = 2'b11;
		14'h0779: color = 2'b11;
		14'h077a: color = 2'b11;
		14'h077b: color = 2'b11;
		14'h077c: color = 2'b11;
		14'h077d: color = 2'b11;
		14'h077e: color = 2'b11;
		14'h077f: color = 2'b11;
		14'h0780: color = 2'b11;
		14'h0781: color = 2'b11;
		14'h0782: color = 2'b11;
		14'h0783: color = 2'b11;
		14'h0784: color = 2'b11;
		14'h0785: color = 2'b11;
		14'h0786: color = 2'b11;
		14'h0787: color = 2'b11;
		14'h0788: color = 2'b11;
		14'h0789: color = 2'b11;
		14'h078a: color = 2'b11;
		14'h078b: color = 2'b11;
		14'h078c: color = 2'b11;
		14'h078d: color = 2'b11;
		14'h078e: color = 2'b11;
		14'h078f: color = 2'b11;
		14'h0790: color = 2'b11;
		14'h0791: color = 2'b11;
		14'h0792: color = 2'b11;
		14'h0793: color = 2'b11;
		14'h0794: color = 2'b11;
		14'h0795: color = 2'b11;
		14'h0796: color = 2'b11;
		14'h0797: color = 2'b11;
		14'h0798: color = 2'b11;
		14'h0799: color = 2'b11;
		14'h079a: color = 2'b11;
		14'h079b: color = 2'b11;
		14'h079c: color = 2'b11;
		14'h079d: color = 2'b11;
		14'h079e: color = 2'b11;
		14'h079f: color = 2'b11;
		14'h07a0: color = 2'b11;
		14'h07a1: color = 2'b11;
		14'h07a2: color = 2'b11;
		14'h07a3: color = 2'b11;
		14'h07a4: color = 2'b11;
		14'h07a5: color = 2'b11;
		14'h07a6: color = 2'b11;
		14'h07a7: color = 2'b11;
		14'h07a8: color = 2'b11;
		14'h07a9: color = 2'b11;
		14'h07aa: color = 2'b11;
		14'h07ab: color = 2'b11;
		14'h07ac: color = 2'b00;
		14'h07ad: color = 2'b00;
		14'h07ae: color = 2'b00;
		14'h07af: color = 2'b00;
		14'h07b0: color = 2'b01;
		14'h07b1: color = 2'b00;
		14'h07b2: color = 2'b00;
		14'h07b3: color = 2'b00;
		14'h07b4: color = 2'b01;
		14'h07b5: color = 2'b00;
		14'h07b6: color = 2'b01;
		14'h07b7: color = 2'b00;
		14'h07b8: color = 2'b00;
		14'h07b9: color = 2'b00;
		14'h07ba: color = 2'b00;
		14'h07bb: color = 2'b00;
		14'h07bc: color = 2'b00;
		14'h07bd: color = 2'b00;
		14'h07be: color = 2'b00;
		14'h07bf: color = 2'b00;
		14'h07c0: color = 2'b00;
		14'h07c1: color = 2'b00;
		14'h07c2: color = 2'b00;
		14'h07c3: color = 2'b00;
		14'h07c4: color = 2'b00;
		14'h07c5: color = 2'b00;
		14'h07c6: color = 2'b00;
		14'h07c7: color = 2'b00;
		14'h07c8: color = 2'b00;
		14'h07c9: color = 2'b00;
		14'h07ca: color = 2'b00;
		14'h07cb: color = 2'b00;
		14'h07cc: color = 2'b00;
		14'h07cd: color = 2'b00;
		14'h07ce: color = 2'b00;
		14'h07cf: color = 2'b00;
		14'h07d0: color = 2'b00;
		14'h07d1: color = 2'b00;
		14'h07d2: color = 2'b00;
		14'h07d3: color = 2'b01;
		14'h07d4: color = 2'b00;
		14'h07d5: color = 2'b00;
		14'h07d6: color = 2'b00;
		14'h07d7: color = 2'b00;
		14'h07d8: color = 2'b00;
		14'h07d9: color = 2'b00;
		14'h07da: color = 2'b00;
		14'h07db: color = 2'b00;
		14'h07dc: color = 2'b00;
		14'h07dd: color = 2'b00;
		14'h07de: color = 2'b00;
		14'h07df: color = 2'b00;
		14'h07e0: color = 2'b00;
		14'h07e1: color = 2'b10;
		14'h07e2: color = 2'b11;
		14'h07e3: color = 2'b11;
		14'h07e4: color = 2'b11;
		14'h07e5: color = 2'b11;
		14'h07e6: color = 2'b11;
		14'h07e7: color = 2'b11;
		14'h07e8: color = 2'b11;
		14'h07e9: color = 2'b11;
		14'h07ea: color = 2'b11;
		14'h07eb: color = 2'b11;
		14'h07ec: color = 2'b11;
		14'h07ed: color = 2'b11;
		14'h07ee: color = 2'b11;
		14'h07ef: color = 2'b11;
		14'h07f0: color = 2'b11;
		14'h07f1: color = 2'b11;
		14'h07f2: color = 2'b11;
		14'h07f3: color = 2'b11;
		14'h07f4: color = 2'b11;
		14'h07f5: color = 2'b11;
		14'h07f6: color = 2'b11;
		14'h07f7: color = 2'b11;
		14'h07f8: color = 2'b11;
		14'h07f9: color = 2'b11;
		14'h07fa: color = 2'b11;
		14'h07fb: color = 2'b11;
		14'h07fc: color = 2'b11;
		14'h07fd: color = 2'b11;
		14'h07fe: color = 2'b11;
		14'h07ff: color = 2'b11;
		14'h0800: color = 2'b11;
		14'h0801: color = 2'b11;
		14'h0802: color = 2'b11;
		14'h0803: color = 2'b11;
		14'h0804: color = 2'b11;
		14'h0805: color = 2'b11;
		14'h0806: color = 2'b11;
		14'h0807: color = 2'b11;
		14'h0808: color = 2'b11;
		14'h0809: color = 2'b11;
		14'h080a: color = 2'b11;
		14'h080b: color = 2'b11;
		14'h080c: color = 2'b11;
		14'h080d: color = 2'b11;
		14'h080e: color = 2'b11;
		14'h080f: color = 2'b11;
		14'h0810: color = 2'b11;
		14'h0811: color = 2'b11;
		14'h0812: color = 2'b11;
		14'h0813: color = 2'b11;
		14'h0814: color = 2'b11;
		14'h0815: color = 2'b11;
		14'h0816: color = 2'b11;
		14'h0817: color = 2'b11;
		14'h0818: color = 2'b11;
		14'h0819: color = 2'b11;
		14'h081a: color = 2'b11;
		14'h081b: color = 2'b11;
		14'h081c: color = 2'b11;
		14'h081d: color = 2'b11;
		14'h081e: color = 2'b11;
		14'h081f: color = 2'b11;
		14'h0820: color = 2'b11;
		14'h0821: color = 2'b11;
		14'h0822: color = 2'b11;
		14'h0823: color = 2'b11;
		14'h0824: color = 2'b11;
		14'h0825: color = 2'b11;
		14'h0826: color = 2'b11;
		14'h0827: color = 2'b11;
		14'h0828: color = 2'b11;
		14'h0829: color = 2'b11;
		14'h082a: color = 2'b11;
		14'h082b: color = 2'b00;
		14'h082c: color = 2'b00;
		14'h082d: color = 2'b00;
		14'h082e: color = 2'b00;
		14'h082f: color = 2'b01;
		14'h0830: color = 2'b00;
		14'h0831: color = 2'b01;
		14'h0832: color = 2'b01;
		14'h0833: color = 2'b01;
		14'h0834: color = 2'b01;
		14'h0835: color = 2'b00;
		14'h0836: color = 2'b00;
		14'h0837: color = 2'b00;
		14'h0838: color = 2'b00;
		14'h0839: color = 2'b00;
		14'h083a: color = 2'b00;
		14'h083b: color = 2'b00;
		14'h083c: color = 2'b00;
		14'h083d: color = 2'b00;
		14'h083e: color = 2'b01;
		14'h083f: color = 2'b00;
		14'h0840: color = 2'b01;
		14'h0841: color = 2'b00;
		14'h0842: color = 2'b00;
		14'h0843: color = 2'b01;
		14'h0844: color = 2'b00;
		14'h0845: color = 2'b00;
		14'h0846: color = 2'b00;
		14'h0847: color = 2'b00;
		14'h0848: color = 2'b00;
		14'h0849: color = 2'b00;
		14'h084a: color = 2'b00;
		14'h084b: color = 2'b00;
		14'h084c: color = 2'b00;
		14'h084d: color = 2'b00;
		14'h084e: color = 2'b00;
		14'h084f: color = 2'b00;
		14'h0850: color = 2'b00;
		14'h0851: color = 2'b00;
		14'h0852: color = 2'b00;
		14'h0853: color = 2'b00;
		14'h0854: color = 2'b01;
		14'h0855: color = 2'b00;
		14'h0856: color = 2'b00;
		14'h0857: color = 2'b00;
		14'h0858: color = 2'b00;
		14'h0859: color = 2'b00;
		14'h085a: color = 2'b00;
		14'h085b: color = 2'b00;
		14'h085c: color = 2'b00;
		14'h085d: color = 2'b00;
		14'h085e: color = 2'b00;
		14'h085f: color = 2'b00;
		14'h0860: color = 2'b00;
		14'h0861: color = 2'b00;
		14'h0862: color = 2'b11;
		14'h0863: color = 2'b11;
		14'h0864: color = 2'b11;
		14'h0865: color = 2'b11;
		14'h0866: color = 2'b11;
		14'h0867: color = 2'b11;
		14'h0868: color = 2'b11;
		14'h0869: color = 2'b11;
		14'h086a: color = 2'b11;
		14'h086b: color = 2'b11;
		14'h086c: color = 2'b11;
		14'h086d: color = 2'b11;
		14'h086e: color = 2'b11;
		14'h086f: color = 2'b11;
		14'h0870: color = 2'b11;
		14'h0871: color = 2'b11;
		14'h0872: color = 2'b11;
		14'h0873: color = 2'b11;
		14'h0874: color = 2'b11;
		14'h0875: color = 2'b11;
		14'h0876: color = 2'b11;
		14'h0877: color = 2'b11;
		14'h0878: color = 2'b11;
		14'h0879: color = 2'b11;
		14'h087a: color = 2'b11;
		14'h087b: color = 2'b11;
		14'h087c: color = 2'b11;
		14'h087d: color = 2'b11;
		14'h087e: color = 2'b11;
		14'h087f: color = 2'b11;
		14'h0880: color = 2'b11;
		14'h0881: color = 2'b11;
		14'h0882: color = 2'b11;
		14'h0883: color = 2'b11;
		14'h0884: color = 2'b11;
		14'h0885: color = 2'b11;
		14'h0886: color = 2'b11;
		14'h0887: color = 2'b11;
		14'h0888: color = 2'b11;
		14'h0889: color = 2'b11;
		14'h088a: color = 2'b11;
		14'h088b: color = 2'b11;
		14'h088c: color = 2'b11;
		14'h088d: color = 2'b11;
		14'h088e: color = 2'b11;
		14'h088f: color = 2'b11;
		14'h0890: color = 2'b11;
		14'h0891: color = 2'b11;
		14'h0892: color = 2'b11;
		14'h0893: color = 2'b11;
		14'h0894: color = 2'b11;
		14'h0895: color = 2'b11;
		14'h0896: color = 2'b11;
		14'h0897: color = 2'b11;
		14'h0898: color = 2'b11;
		14'h0899: color = 2'b11;
		14'h089a: color = 2'b11;
		14'h089b: color = 2'b11;
		14'h089c: color = 2'b11;
		14'h089d: color = 2'b11;
		14'h089e: color = 2'b11;
		14'h089f: color = 2'b11;
		14'h08a0: color = 2'b11;
		14'h08a1: color = 2'b11;
		14'h08a2: color = 2'b11;
		14'h08a3: color = 2'b11;
		14'h08a4: color = 2'b11;
		14'h08a5: color = 2'b11;
		14'h08a6: color = 2'b11;
		14'h08a7: color = 2'b11;
		14'h08a8: color = 2'b11;
		14'h08a9: color = 2'b11;
		14'h08aa: color = 2'b00;
		14'h08ab: color = 2'b00;
		14'h08ac: color = 2'b00;
		14'h08ad: color = 2'b01;
		14'h08ae: color = 2'b00;
		14'h08af: color = 2'b00;
		14'h08b0: color = 2'b01;
		14'h08b1: color = 2'b00;
		14'h08b2: color = 2'b01;
		14'h08b3: color = 2'b00;
		14'h08b4: color = 2'b01;
		14'h08b5: color = 2'b01;
		14'h08b6: color = 2'b00;
		14'h08b7: color = 2'b00;
		14'h08b8: color = 2'b00;
		14'h08b9: color = 2'b00;
		14'h08ba: color = 2'b01;
		14'h08bb: color = 2'b00;
		14'h08bc: color = 2'b01;
		14'h08bd: color = 2'b01;
		14'h08be: color = 2'b00;
		14'h08bf: color = 2'b01;
		14'h08c0: color = 2'b00;
		14'h08c1: color = 2'b00;
		14'h08c2: color = 2'b00;
		14'h08c3: color = 2'b00;
		14'h08c4: color = 2'b00;
		14'h08c5: color = 2'b00;
		14'h08c6: color = 2'b00;
		14'h08c7: color = 2'b00;
		14'h08c8: color = 2'b00;
		14'h08c9: color = 2'b00;
		14'h08ca: color = 2'b00;
		14'h08cb: color = 2'b00;
		14'h08cc: color = 2'b00;
		14'h08cd: color = 2'b00;
		14'h08ce: color = 2'b00;
		14'h08cf: color = 2'b00;
		14'h08d0: color = 2'b00;
		14'h08d1: color = 2'b00;
		14'h08d2: color = 2'b00;
		14'h08d3: color = 2'b00;
		14'h08d4: color = 2'b00;
		14'h08d5: color = 2'b00;
		14'h08d6: color = 2'b00;
		14'h08d7: color = 2'b00;
		14'h08d8: color = 2'b00;
		14'h08d9: color = 2'b00;
		14'h08da: color = 2'b00;
		14'h08db: color = 2'b00;
		14'h08dc: color = 2'b00;
		14'h08dd: color = 2'b00;
		14'h08de: color = 2'b00;
		14'h08df: color = 2'b00;
		14'h08e0: color = 2'b00;
		14'h08e1: color = 2'b00;
		14'h08e2: color = 2'b10;
		14'h08e3: color = 2'b11;
		14'h08e4: color = 2'b11;
		14'h08e5: color = 2'b11;
		14'h08e6: color = 2'b11;
		14'h08e7: color = 2'b11;
		14'h08e8: color = 2'b11;
		14'h08e9: color = 2'b11;
		14'h08ea: color = 2'b11;
		14'h08eb: color = 2'b11;
		14'h08ec: color = 2'b11;
		14'h08ed: color = 2'b11;
		14'h08ee: color = 2'b11;
		14'h08ef: color = 2'b11;
		14'h08f0: color = 2'b11;
		14'h08f1: color = 2'b11;
		14'h08f2: color = 2'b11;
		14'h08f3: color = 2'b11;
		14'h08f4: color = 2'b11;
		14'h08f5: color = 2'b11;
		14'h08f6: color = 2'b11;
		14'h08f7: color = 2'b11;
		14'h08f8: color = 2'b11;
		14'h08f9: color = 2'b11;
		14'h08fa: color = 2'b11;
		14'h08fb: color = 2'b11;
		14'h08fc: color = 2'b11;
		14'h08fd: color = 2'b11;
		14'h08fe: color = 2'b11;
		14'h08ff: color = 2'b11;
		14'h0900: color = 2'b11;
		14'h0901: color = 2'b11;
		14'h0902: color = 2'b11;
		14'h0903: color = 2'b11;
		14'h0904: color = 2'b11;
		14'h0905: color = 2'b11;
		14'h0906: color = 2'b11;
		14'h0907: color = 2'b11;
		14'h0908: color = 2'b11;
		14'h0909: color = 2'b11;
		14'h090a: color = 2'b11;
		14'h090b: color = 2'b11;
		14'h090c: color = 2'b11;
		14'h090d: color = 2'b11;
		14'h090e: color = 2'b11;
		14'h090f: color = 2'b11;
		14'h0910: color = 2'b11;
		14'h0911: color = 2'b11;
		14'h0912: color = 2'b11;
		14'h0913: color = 2'b11;
		14'h0914: color = 2'b11;
		14'h0915: color = 2'b11;
		14'h0916: color = 2'b11;
		14'h0917: color = 2'b11;
		14'h0918: color = 2'b11;
		14'h0919: color = 2'b11;
		14'h091a: color = 2'b11;
		14'h091b: color = 2'b11;
		14'h091c: color = 2'b11;
		14'h091d: color = 2'b11;
		14'h091e: color = 2'b11;
		14'h091f: color = 2'b11;
		14'h0920: color = 2'b11;
		14'h0921: color = 2'b11;
		14'h0922: color = 2'b11;
		14'h0923: color = 2'b11;
		14'h0924: color = 2'b11;
		14'h0925: color = 2'b11;
		14'h0926: color = 2'b11;
		14'h0927: color = 2'b11;
		14'h0928: color = 2'b11;
		14'h0929: color = 2'b10;
		14'h092a: color = 2'b00;
		14'h092b: color = 2'b00;
		14'h092c: color = 2'b00;
		14'h092d: color = 2'b01;
		14'h092e: color = 2'b00;
		14'h092f: color = 2'b01;
		14'h0930: color = 2'b00;
		14'h0931: color = 2'b01;
		14'h0932: color = 2'b01;
		14'h0933: color = 2'b00;
		14'h0934: color = 2'b00;
		14'h0935: color = 2'b00;
		14'h0936: color = 2'b00;
		14'h0937: color = 2'b01;
		14'h0938: color = 2'b01;
		14'h0939: color = 2'b01;
		14'h093a: color = 2'b00;
		14'h093b: color = 2'b01;
		14'h093c: color = 2'b00;
		14'h093d: color = 2'b00;
		14'h093e: color = 2'b01;
		14'h093f: color = 2'b00;
		14'h0940: color = 2'b00;
		14'h0941: color = 2'b01;
		14'h0942: color = 2'b00;
		14'h0943: color = 2'b00;
		14'h0944: color = 2'b00;
		14'h0945: color = 2'b00;
		14'h0946: color = 2'b00;
		14'h0947: color = 2'b00;
		14'h0948: color = 2'b00;
		14'h0949: color = 2'b00;
		14'h094a: color = 2'b00;
		14'h094b: color = 2'b00;
		14'h094c: color = 2'b00;
		14'h094d: color = 2'b00;
		14'h094e: color = 2'b00;
		14'h094f: color = 2'b00;
		14'h0950: color = 2'b00;
		14'h0951: color = 2'b00;
		14'h0952: color = 2'b00;
		14'h0953: color = 2'b00;
		14'h0954: color = 2'b00;
		14'h0955: color = 2'b00;
		14'h0956: color = 2'b00;
		14'h0957: color = 2'b00;
		14'h0958: color = 2'b00;
		14'h0959: color = 2'b00;
		14'h095a: color = 2'b00;
		14'h095b: color = 2'b00;
		14'h095c: color = 2'b00;
		14'h095d: color = 2'b00;
		14'h095e: color = 2'b00;
		14'h095f: color = 2'b00;
		14'h0960: color = 2'b00;
		14'h0961: color = 2'b00;
		14'h0962: color = 2'b00;
		14'h0963: color = 2'b11;
		14'h0964: color = 2'b11;
		14'h0965: color = 2'b11;
		14'h0966: color = 2'b11;
		14'h0967: color = 2'b11;
		14'h0968: color = 2'b11;
		14'h0969: color = 2'b11;
		14'h096a: color = 2'b11;
		14'h096b: color = 2'b11;
		14'h096c: color = 2'b11;
		14'h096d: color = 2'b11;
		14'h096e: color = 2'b11;
		14'h096f: color = 2'b11;
		14'h0970: color = 2'b11;
		14'h0971: color = 2'b11;
		14'h0972: color = 2'b11;
		14'h0973: color = 2'b11;
		14'h0974: color = 2'b11;
		14'h0975: color = 2'b11;
		14'h0976: color = 2'b11;
		14'h0977: color = 2'b11;
		14'h0978: color = 2'b11;
		14'h0979: color = 2'b11;
		14'h097a: color = 2'b11;
		14'h097b: color = 2'b11;
		14'h097c: color = 2'b11;
		14'h097d: color = 2'b11;
		14'h097e: color = 2'b11;
		14'h097f: color = 2'b11;
		14'h0980: color = 2'b11;
		14'h0981: color = 2'b11;
		14'h0982: color = 2'b11;
		14'h0983: color = 2'b11;
		14'h0984: color = 2'b11;
		14'h0985: color = 2'b11;
		14'h0986: color = 2'b11;
		14'h0987: color = 2'b11;
		14'h0988: color = 2'b11;
		14'h0989: color = 2'b11;
		14'h098a: color = 2'b11;
		14'h098b: color = 2'b11;
		14'h098c: color = 2'b11;
		14'h098d: color = 2'b11;
		14'h098e: color = 2'b11;
		14'h098f: color = 2'b11;
		14'h0990: color = 2'b11;
		14'h0991: color = 2'b11;
		14'h0992: color = 2'b11;
		14'h0993: color = 2'b11;
		14'h0994: color = 2'b11;
		14'h0995: color = 2'b11;
		14'h0996: color = 2'b11;
		14'h0997: color = 2'b11;
		14'h0998: color = 2'b11;
		14'h0999: color = 2'b11;
		14'h099a: color = 2'b11;
		14'h099b: color = 2'b11;
		14'h099c: color = 2'b11;
		14'h099d: color = 2'b11;
		14'h099e: color = 2'b11;
		14'h099f: color = 2'b11;
		14'h09a0: color = 2'b11;
		14'h09a1: color = 2'b11;
		14'h09a2: color = 2'b11;
		14'h09a3: color = 2'b11;
		14'h09a4: color = 2'b11;
		14'h09a5: color = 2'b11;
		14'h09a6: color = 2'b11;
		14'h09a7: color = 2'b11;
		14'h09a8: color = 2'b11;
		14'h09a9: color = 2'b01;
		14'h09aa: color = 2'b00;
		14'h09ab: color = 2'b00;
		14'h09ac: color = 2'b00;
		14'h09ad: color = 2'b01;
		14'h09ae: color = 2'b01;
		14'h09af: color = 2'b00;
		14'h09b0: color = 2'b01;
		14'h09b1: color = 2'b01;
		14'h09b2: color = 2'b00;
		14'h09b3: color = 2'b01;
		14'h09b4: color = 2'b00;
		14'h09b5: color = 2'b00;
		14'h09b6: color = 2'b00;
		14'h09b7: color = 2'b01;
		14'h09b8: color = 2'b01;
		14'h09b9: color = 2'b01;
		14'h09ba: color = 2'b01;
		14'h09bb: color = 2'b00;
		14'h09bc: color = 2'b00;
		14'h09bd: color = 2'b01;
		14'h09be: color = 2'b00;
		14'h09bf: color = 2'b00;
		14'h09c0: color = 2'b01;
		14'h09c1: color = 2'b00;
		14'h09c2: color = 2'b01;
		14'h09c3: color = 2'b00;
		14'h09c4: color = 2'b00;
		14'h09c5: color = 2'b00;
		14'h09c6: color = 2'b00;
		14'h09c7: color = 2'b00;
		14'h09c8: color = 2'b00;
		14'h09c9: color = 2'b00;
		14'h09ca: color = 2'b00;
		14'h09cb: color = 2'b00;
		14'h09cc: color = 2'b00;
		14'h09cd: color = 2'b00;
		14'h09ce: color = 2'b00;
		14'h09cf: color = 2'b00;
		14'h09d0: color = 2'b00;
		14'h09d1: color = 2'b00;
		14'h09d2: color = 2'b00;
		14'h09d3: color = 2'b00;
		14'h09d4: color = 2'b00;
		14'h09d5: color = 2'b00;
		14'h09d6: color = 2'b00;
		14'h09d7: color = 2'b00;
		14'h09d8: color = 2'b00;
		14'h09d9: color = 2'b00;
		14'h09da: color = 2'b00;
		14'h09db: color = 2'b00;
		14'h09dc: color = 2'b00;
		14'h09dd: color = 2'b00;
		14'h09de: color = 2'b00;
		14'h09df: color = 2'b00;
		14'h09e0: color = 2'b00;
		14'h09e1: color = 2'b00;
		14'h09e2: color = 2'b00;
		14'h09e3: color = 2'b11;
		14'h09e4: color = 2'b11;
		14'h09e5: color = 2'b11;
		14'h09e6: color = 2'b11;
		14'h09e7: color = 2'b11;
		14'h09e8: color = 2'b11;
		14'h09e9: color = 2'b11;
		14'h09ea: color = 2'b11;
		14'h09eb: color = 2'b11;
		14'h09ec: color = 2'b11;
		14'h09ed: color = 2'b11;
		14'h09ee: color = 2'b11;
		14'h09ef: color = 2'b11;
		14'h09f0: color = 2'b11;
		14'h09f1: color = 2'b11;
		14'h09f2: color = 2'b11;
		14'h09f3: color = 2'b11;
		14'h09f4: color = 2'b11;
		14'h09f5: color = 2'b11;
		14'h09f6: color = 2'b11;
		14'h09f7: color = 2'b11;
		14'h09f8: color = 2'b11;
		14'h09f9: color = 2'b11;
		14'h09fa: color = 2'b11;
		14'h09fb: color = 2'b11;
		14'h09fc: color = 2'b11;
		14'h09fd: color = 2'b11;
		14'h09fe: color = 2'b11;
		14'h09ff: color = 2'b11;
		14'h0a00: color = 2'b11;
		14'h0a01: color = 2'b11;
		14'h0a02: color = 2'b11;
		14'h0a03: color = 2'b11;
		14'h0a04: color = 2'b11;
		14'h0a05: color = 2'b11;
		14'h0a06: color = 2'b11;
		14'h0a07: color = 2'b11;
		14'h0a08: color = 2'b11;
		14'h0a09: color = 2'b11;
		14'h0a0a: color = 2'b11;
		14'h0a0b: color = 2'b11;
		14'h0a0c: color = 2'b11;
		14'h0a0d: color = 2'b11;
		14'h0a0e: color = 2'b11;
		14'h0a0f: color = 2'b11;
		14'h0a10: color = 2'b11;
		14'h0a11: color = 2'b11;
		14'h0a12: color = 2'b11;
		14'h0a13: color = 2'b11;
		14'h0a14: color = 2'b11;
		14'h0a15: color = 2'b11;
		14'h0a16: color = 2'b11;
		14'h0a17: color = 2'b11;
		14'h0a18: color = 2'b11;
		14'h0a19: color = 2'b11;
		14'h0a1a: color = 2'b11;
		14'h0a1b: color = 2'b11;
		14'h0a1c: color = 2'b11;
		14'h0a1d: color = 2'b11;
		14'h0a1e: color = 2'b11;
		14'h0a1f: color = 2'b11;
		14'h0a20: color = 2'b11;
		14'h0a21: color = 2'b11;
		14'h0a22: color = 2'b11;
		14'h0a23: color = 2'b11;
		14'h0a24: color = 2'b11;
		14'h0a25: color = 2'b11;
		14'h0a26: color = 2'b11;
		14'h0a27: color = 2'b11;
		14'h0a28: color = 2'b11;
		14'h0a29: color = 2'b01;
		14'h0a2a: color = 2'b00;
		14'h0a2b: color = 2'b00;
		14'h0a2c: color = 2'b01;
		14'h0a2d: color = 2'b01;
		14'h0a2e: color = 2'b00;
		14'h0a2f: color = 2'b00;
		14'h0a30: color = 2'b01;
		14'h0a31: color = 2'b01;
		14'h0a32: color = 2'b01;
		14'h0a33: color = 2'b00;
		14'h0a34: color = 2'b00;
		14'h0a35: color = 2'b01;
		14'h0a36: color = 2'b01;
		14'h0a37: color = 2'b01;
		14'h0a38: color = 2'b01;
		14'h0a39: color = 2'b01;
		14'h0a3a: color = 2'b00;
		14'h0a3b: color = 2'b00;
		14'h0a3c: color = 2'b01;
		14'h0a3d: color = 2'b00;
		14'h0a3e: color = 2'b00;
		14'h0a3f: color = 2'b00;
		14'h0a40: color = 2'b00;
		14'h0a41: color = 2'b00;
		14'h0a42: color = 2'b01;
		14'h0a43: color = 2'b00;
		14'h0a44: color = 2'b00;
		14'h0a45: color = 2'b00;
		14'h0a46: color = 2'b00;
		14'h0a47: color = 2'b00;
		14'h0a48: color = 2'b00;
		14'h0a49: color = 2'b00;
		14'h0a4a: color = 2'b00;
		14'h0a4b: color = 2'b00;
		14'h0a4c: color = 2'b00;
		14'h0a4d: color = 2'b00;
		14'h0a4e: color = 2'b00;
		14'h0a4f: color = 2'b00;
		14'h0a50: color = 2'b00;
		14'h0a51: color = 2'b00;
		14'h0a52: color = 2'b00;
		14'h0a53: color = 2'b00;
		14'h0a54: color = 2'b00;
		14'h0a55: color = 2'b00;
		14'h0a56: color = 2'b00;
		14'h0a57: color = 2'b00;
		14'h0a58: color = 2'b00;
		14'h0a59: color = 2'b00;
		14'h0a5a: color = 2'b00;
		14'h0a5b: color = 2'b00;
		14'h0a5c: color = 2'b00;
		14'h0a5d: color = 2'b00;
		14'h0a5e: color = 2'b00;
		14'h0a5f: color = 2'b00;
		14'h0a60: color = 2'b00;
		14'h0a61: color = 2'b00;
		14'h0a62: color = 2'b00;
		14'h0a63: color = 2'b00;
		14'h0a64: color = 2'b11;
		14'h0a65: color = 2'b11;
		14'h0a66: color = 2'b11;
		14'h0a67: color = 2'b11;
		14'h0a68: color = 2'b11;
		14'h0a69: color = 2'b11;
		14'h0a6a: color = 2'b11;
		14'h0a6b: color = 2'b11;
		14'h0a6c: color = 2'b11;
		14'h0a6d: color = 2'b11;
		14'h0a6e: color = 2'b11;
		14'h0a6f: color = 2'b11;
		14'h0a70: color = 2'b11;
		14'h0a71: color = 2'b11;
		14'h0a72: color = 2'b11;
		14'h0a73: color = 2'b11;
		14'h0a74: color = 2'b11;
		14'h0a75: color = 2'b11;
		14'h0a76: color = 2'b11;
		14'h0a77: color = 2'b11;
		14'h0a78: color = 2'b11;
		14'h0a79: color = 2'b11;
		14'h0a7a: color = 2'b11;
		14'h0a7b: color = 2'b11;
		14'h0a7c: color = 2'b11;
		14'h0a7d: color = 2'b11;
		14'h0a7e: color = 2'b11;
		14'h0a7f: color = 2'b11;
		14'h0a80: color = 2'b11;
		14'h0a81: color = 2'b11;
		14'h0a82: color = 2'b11;
		14'h0a83: color = 2'b11;
		14'h0a84: color = 2'b11;
		14'h0a85: color = 2'b11;
		14'h0a86: color = 2'b11;
		14'h0a87: color = 2'b11;
		14'h0a88: color = 2'b11;
		14'h0a89: color = 2'b11;
		14'h0a8a: color = 2'b11;
		14'h0a8b: color = 2'b11;
		14'h0a8c: color = 2'b11;
		14'h0a8d: color = 2'b11;
		14'h0a8e: color = 2'b11;
		14'h0a8f: color = 2'b11;
		14'h0a90: color = 2'b11;
		14'h0a91: color = 2'b11;
		14'h0a92: color = 2'b11;
		14'h0a93: color = 2'b11;
		14'h0a94: color = 2'b11;
		14'h0a95: color = 2'b11;
		14'h0a96: color = 2'b11;
		14'h0a97: color = 2'b11;
		14'h0a98: color = 2'b11;
		14'h0a99: color = 2'b11;
		14'h0a9a: color = 2'b11;
		14'h0a9b: color = 2'b11;
		14'h0a9c: color = 2'b11;
		14'h0a9d: color = 2'b11;
		14'h0a9e: color = 2'b11;
		14'h0a9f: color = 2'b11;
		14'h0aa0: color = 2'b11;
		14'h0aa1: color = 2'b11;
		14'h0aa2: color = 2'b11;
		14'h0aa3: color = 2'b11;
		14'h0aa4: color = 2'b11;
		14'h0aa5: color = 2'b11;
		14'h0aa6: color = 2'b11;
		14'h0aa7: color = 2'b11;
		14'h0aa8: color = 2'b11;
		14'h0aa9: color = 2'b00;
		14'h0aaa: color = 2'b00;
		14'h0aab: color = 2'b00;
		14'h0aac: color = 2'b00;
		14'h0aad: color = 2'b01;
		14'h0aae: color = 2'b00;
		14'h0aaf: color = 2'b00;
		14'h0ab0: color = 2'b00;
		14'h0ab1: color = 2'b01;
		14'h0ab2: color = 2'b01;
		14'h0ab3: color = 2'b00;
		14'h0ab4: color = 2'b00;
		14'h0ab5: color = 2'b01;
		14'h0ab6: color = 2'b01;
		14'h0ab7: color = 2'b01;
		14'h0ab8: color = 2'b01;
		14'h0ab9: color = 2'b00;
		14'h0aba: color = 2'b00;
		14'h0abb: color = 2'b00;
		14'h0abc: color = 2'b00;
		14'h0abd: color = 2'b00;
		14'h0abe: color = 2'b00;
		14'h0abf: color = 2'b00;
		14'h0ac0: color = 2'b00;
		14'h0ac1: color = 2'b00;
		14'h0ac2: color = 2'b00;
		14'h0ac3: color = 2'b00;
		14'h0ac4: color = 2'b00;
		14'h0ac5: color = 2'b00;
		14'h0ac6: color = 2'b00;
		14'h0ac7: color = 2'b00;
		14'h0ac8: color = 2'b00;
		14'h0ac9: color = 2'b00;
		14'h0aca: color = 2'b00;
		14'h0acb: color = 2'b00;
		14'h0acc: color = 2'b00;
		14'h0acd: color = 2'b00;
		14'h0ace: color = 2'b00;
		14'h0acf: color = 2'b00;
		14'h0ad0: color = 2'b00;
		14'h0ad1: color = 2'b00;
		14'h0ad2: color = 2'b00;
		14'h0ad3: color = 2'b00;
		14'h0ad4: color = 2'b00;
		14'h0ad5: color = 2'b00;
		14'h0ad6: color = 2'b00;
		14'h0ad7: color = 2'b00;
		14'h0ad8: color = 2'b00;
		14'h0ad9: color = 2'b00;
		14'h0ada: color = 2'b00;
		14'h0adb: color = 2'b00;
		14'h0adc: color = 2'b00;
		14'h0add: color = 2'b00;
		14'h0ade: color = 2'b00;
		14'h0adf: color = 2'b00;
		14'h0ae0: color = 2'b00;
		14'h0ae1: color = 2'b00;
		14'h0ae2: color = 2'b00;
		14'h0ae3: color = 2'b00;
		14'h0ae4: color = 2'b10;
		14'h0ae5: color = 2'b11;
		14'h0ae6: color = 2'b11;
		14'h0ae7: color = 2'b11;
		14'h0ae8: color = 2'b11;
		14'h0ae9: color = 2'b11;
		14'h0aea: color = 2'b11;
		14'h0aeb: color = 2'b11;
		14'h0aec: color = 2'b11;
		14'h0aed: color = 2'b11;
		14'h0aee: color = 2'b11;
		14'h0aef: color = 2'b11;
		14'h0af0: color = 2'b11;
		14'h0af1: color = 2'b11;
		14'h0af2: color = 2'b11;
		14'h0af3: color = 2'b11;
		14'h0af4: color = 2'b11;
		14'h0af5: color = 2'b11;
		14'h0af6: color = 2'b11;
		14'h0af7: color = 2'b11;
		14'h0af8: color = 2'b11;
		14'h0af9: color = 2'b11;
		14'h0afa: color = 2'b11;
		14'h0afb: color = 2'b11;
		14'h0afc: color = 2'b11;
		14'h0afd: color = 2'b11;
		14'h0afe: color = 2'b11;
		14'h0aff: color = 2'b11;
		14'h0b00: color = 2'b11;
		14'h0b01: color = 2'b11;
		14'h0b02: color = 2'b11;
		14'h0b03: color = 2'b11;
		14'h0b04: color = 2'b11;
		14'h0b05: color = 2'b11;
		14'h0b06: color = 2'b11;
		14'h0b07: color = 2'b11;
		14'h0b08: color = 2'b11;
		14'h0b09: color = 2'b11;
		14'h0b0a: color = 2'b11;
		14'h0b0b: color = 2'b11;
		14'h0b0c: color = 2'b11;
		14'h0b0d: color = 2'b11;
		14'h0b0e: color = 2'b11;
		14'h0b0f: color = 2'b11;
		14'h0b10: color = 2'b11;
		14'h0b11: color = 2'b11;
		14'h0b12: color = 2'b11;
		14'h0b13: color = 2'b11;
		14'h0b14: color = 2'b11;
		14'h0b15: color = 2'b11;
		14'h0b16: color = 2'b11;
		14'h0b17: color = 2'b11;
		14'h0b18: color = 2'b11;
		14'h0b19: color = 2'b11;
		14'h0b1a: color = 2'b11;
		14'h0b1b: color = 2'b11;
		14'h0b1c: color = 2'b11;
		14'h0b1d: color = 2'b11;
		14'h0b1e: color = 2'b11;
		14'h0b1f: color = 2'b11;
		14'h0b20: color = 2'b11;
		14'h0b21: color = 2'b11;
		14'h0b22: color = 2'b11;
		14'h0b23: color = 2'b11;
		14'h0b24: color = 2'b11;
		14'h0b25: color = 2'b11;
		14'h0b26: color = 2'b01;
		14'h0b27: color = 2'b00;
		14'h0b28: color = 2'b00;
		14'h0b29: color = 2'b00;
		14'h0b2a: color = 2'b00;
		14'h0b2b: color = 2'b00;
		14'h0b2c: color = 2'b00;
		14'h0b2d: color = 2'b00;
		14'h0b2e: color = 2'b00;
		14'h0b2f: color = 2'b00;
		14'h0b30: color = 2'b00;
		14'h0b31: color = 2'b01;
		14'h0b32: color = 2'b00;
		14'h0b33: color = 2'b01;
		14'h0b34: color = 2'b00;
		14'h0b35: color = 2'b00;
		14'h0b36: color = 2'b00;
		14'h0b37: color = 2'b00;
		14'h0b38: color = 2'b00;
		14'h0b39: color = 2'b00;
		14'h0b3a: color = 2'b00;
		14'h0b3b: color = 2'b00;
		14'h0b3c: color = 2'b00;
		14'h0b3d: color = 2'b00;
		14'h0b3e: color = 2'b00;
		14'h0b3f: color = 2'b00;
		14'h0b40: color = 2'b00;
		14'h0b41: color = 2'b00;
		14'h0b42: color = 2'b00;
		14'h0b43: color = 2'b01;
		14'h0b44: color = 2'b00;
		14'h0b45: color = 2'b00;
		14'h0b46: color = 2'b00;
		14'h0b47: color = 2'b00;
		14'h0b48: color = 2'b00;
		14'h0b49: color = 2'b00;
		14'h0b4a: color = 2'b00;
		14'h0b4b: color = 2'b00;
		14'h0b4c: color = 2'b00;
		14'h0b4d: color = 2'b00;
		14'h0b4e: color = 2'b00;
		14'h0b4f: color = 2'b00;
		14'h0b50: color = 2'b00;
		14'h0b51: color = 2'b00;
		14'h0b52: color = 2'b00;
		14'h0b53: color = 2'b00;
		14'h0b54: color = 2'b00;
		14'h0b55: color = 2'b00;
		14'h0b56: color = 2'b00;
		14'h0b57: color = 2'b00;
		14'h0b58: color = 2'b00;
		14'h0b59: color = 2'b00;
		14'h0b5a: color = 2'b00;
		14'h0b5b: color = 2'b00;
		14'h0b5c: color = 2'b00;
		14'h0b5d: color = 2'b00;
		14'h0b5e: color = 2'b00;
		14'h0b5f: color = 2'b00;
		14'h0b60: color = 2'b00;
		14'h0b61: color = 2'b00;
		14'h0b62: color = 2'b00;
		14'h0b63: color = 2'b00;
		14'h0b64: color = 2'b10;
		14'h0b65: color = 2'b11;
		14'h0b66: color = 2'b11;
		14'h0b67: color = 2'b11;
		14'h0b68: color = 2'b11;
		14'h0b69: color = 2'b11;
		14'h0b6a: color = 2'b11;
		14'h0b6b: color = 2'b11;
		14'h0b6c: color = 2'b11;
		14'h0b6d: color = 2'b11;
		14'h0b6e: color = 2'b11;
		14'h0b6f: color = 2'b11;
		14'h0b70: color = 2'b11;
		14'h0b71: color = 2'b11;
		14'h0b72: color = 2'b11;
		14'h0b73: color = 2'b11;
		14'h0b74: color = 2'b11;
		14'h0b75: color = 2'b11;
		14'h0b76: color = 2'b11;
		14'h0b77: color = 2'b11;
		14'h0b78: color = 2'b11;
		14'h0b79: color = 2'b11;
		14'h0b7a: color = 2'b11;
		14'h0b7b: color = 2'b11;
		14'h0b7c: color = 2'b11;
		14'h0b7d: color = 2'b11;
		14'h0b7e: color = 2'b11;
		14'h0b7f: color = 2'b11;
		14'h0b80: color = 2'b11;
		14'h0b81: color = 2'b11;
		14'h0b82: color = 2'b11;
		14'h0b83: color = 2'b11;
		14'h0b84: color = 2'b11;
		14'h0b85: color = 2'b11;
		14'h0b86: color = 2'b11;
		14'h0b87: color = 2'b11;
		14'h0b88: color = 2'b11;
		14'h0b89: color = 2'b11;
		14'h0b8a: color = 2'b11;
		14'h0b8b: color = 2'b11;
		14'h0b8c: color = 2'b11;
		14'h0b8d: color = 2'b11;
		14'h0b8e: color = 2'b11;
		14'h0b8f: color = 2'b11;
		14'h0b90: color = 2'b11;
		14'h0b91: color = 2'b11;
		14'h0b92: color = 2'b11;
		14'h0b93: color = 2'b11;
		14'h0b94: color = 2'b11;
		14'h0b95: color = 2'b11;
		14'h0b96: color = 2'b11;
		14'h0b97: color = 2'b11;
		14'h0b98: color = 2'b11;
		14'h0b99: color = 2'b11;
		14'h0b9a: color = 2'b11;
		14'h0b9b: color = 2'b11;
		14'h0b9c: color = 2'b11;
		14'h0b9d: color = 2'b11;
		14'h0b9e: color = 2'b11;
		14'h0b9f: color = 2'b11;
		14'h0ba0: color = 2'b11;
		14'h0ba1: color = 2'b11;
		14'h0ba2: color = 2'b11;
		14'h0ba3: color = 2'b11;
		14'h0ba4: color = 2'b11;
		14'h0ba5: color = 2'b11;
		14'h0ba6: color = 2'b01;
		14'h0ba7: color = 2'b00;
		14'h0ba8: color = 2'b00;
		14'h0ba9: color = 2'b00;
		14'h0baa: color = 2'b00;
		14'h0bab: color = 2'b00;
		14'h0bac: color = 2'b00;
		14'h0bad: color = 2'b00;
		14'h0bae: color = 2'b01;
		14'h0baf: color = 2'b00;
		14'h0bb0: color = 2'b00;
		14'h0bb1: color = 2'b00;
		14'h0bb2: color = 2'b00;
		14'h0bb3: color = 2'b01;
		14'h0bb4: color = 2'b00;
		14'h0bb5: color = 2'b01;
		14'h0bb6: color = 2'b00;
		14'h0bb7: color = 2'b00;
		14'h0bb8: color = 2'b00;
		14'h0bb9: color = 2'b00;
		14'h0bba: color = 2'b00;
		14'h0bbb: color = 2'b00;
		14'h0bbc: color = 2'b00;
		14'h0bbd: color = 2'b00;
		14'h0bbe: color = 2'b00;
		14'h0bbf: color = 2'b00;
		14'h0bc0: color = 2'b00;
		14'h0bc1: color = 2'b00;
		14'h0bc2: color = 2'b00;
		14'h0bc3: color = 2'b00;
		14'h0bc4: color = 2'b00;
		14'h0bc5: color = 2'b00;
		14'h0bc6: color = 2'b00;
		14'h0bc7: color = 2'b00;
		14'h0bc8: color = 2'b00;
		14'h0bc9: color = 2'b00;
		14'h0bca: color = 2'b00;
		14'h0bcb: color = 2'b00;
		14'h0bcc: color = 2'b00;
		14'h0bcd: color = 2'b00;
		14'h0bce: color = 2'b00;
		14'h0bcf: color = 2'b00;
		14'h0bd0: color = 2'b00;
		14'h0bd1: color = 2'b00;
		14'h0bd2: color = 2'b00;
		14'h0bd3: color = 2'b00;
		14'h0bd4: color = 2'b00;
		14'h0bd5: color = 2'b00;
		14'h0bd6: color = 2'b00;
		14'h0bd7: color = 2'b00;
		14'h0bd8: color = 2'b00;
		14'h0bd9: color = 2'b00;
		14'h0bda: color = 2'b00;
		14'h0bdb: color = 2'b00;
		14'h0bdc: color = 2'b00;
		14'h0bdd: color = 2'b00;
		14'h0bde: color = 2'b00;
		14'h0bdf: color = 2'b00;
		14'h0be0: color = 2'b00;
		14'h0be1: color = 2'b00;
		14'h0be2: color = 2'b00;
		14'h0be3: color = 2'b00;
		14'h0be4: color = 2'b00;
		14'h0be5: color = 2'b11;
		14'h0be6: color = 2'b11;
		14'h0be7: color = 2'b11;
		14'h0be8: color = 2'b11;
		14'h0be9: color = 2'b11;
		14'h0bea: color = 2'b11;
		14'h0beb: color = 2'b11;
		14'h0bec: color = 2'b11;
		14'h0bed: color = 2'b11;
		14'h0bee: color = 2'b11;
		14'h0bef: color = 2'b11;
		14'h0bf0: color = 2'b11;
		14'h0bf1: color = 2'b11;
		14'h0bf2: color = 2'b11;
		14'h0bf3: color = 2'b11;
		14'h0bf4: color = 2'b11;
		14'h0bf5: color = 2'b11;
		14'h0bf6: color = 2'b11;
		14'h0bf7: color = 2'b11;
		14'h0bf8: color = 2'b11;
		14'h0bf9: color = 2'b11;
		14'h0bfa: color = 2'b11;
		14'h0bfb: color = 2'b11;
		14'h0bfc: color = 2'b11;
		14'h0bfd: color = 2'b11;
		14'h0bfe: color = 2'b11;
		14'h0bff: color = 2'b11;
		14'h0c00: color = 2'b11;
		14'h0c01: color = 2'b11;
		14'h0c02: color = 2'b11;
		14'h0c03: color = 2'b11;
		14'h0c04: color = 2'b11;
		14'h0c05: color = 2'b11;
		14'h0c06: color = 2'b11;
		14'h0c07: color = 2'b11;
		14'h0c08: color = 2'b11;
		14'h0c09: color = 2'b11;
		14'h0c0a: color = 2'b11;
		14'h0c0b: color = 2'b11;
		14'h0c0c: color = 2'b11;
		14'h0c0d: color = 2'b11;
		14'h0c0e: color = 2'b11;
		14'h0c0f: color = 2'b11;
		14'h0c10: color = 2'b11;
		14'h0c11: color = 2'b11;
		14'h0c12: color = 2'b11;
		14'h0c13: color = 2'b11;
		14'h0c14: color = 2'b11;
		14'h0c15: color = 2'b11;
		14'h0c16: color = 2'b11;
		14'h0c17: color = 2'b11;
		14'h0c18: color = 2'b11;
		14'h0c19: color = 2'b11;
		14'h0c1a: color = 2'b11;
		14'h0c1b: color = 2'b11;
		14'h0c1c: color = 2'b11;
		14'h0c1d: color = 2'b11;
		14'h0c1e: color = 2'b11;
		14'h0c1f: color = 2'b11;
		14'h0c20: color = 2'b11;
		14'h0c21: color = 2'b11;
		14'h0c22: color = 2'b11;
		14'h0c23: color = 2'b11;
		14'h0c24: color = 2'b11;
		14'h0c25: color = 2'b11;
		14'h0c26: color = 2'b01;
		14'h0c27: color = 2'b00;
		14'h0c28: color = 2'b00;
		14'h0c29: color = 2'b00;
		14'h0c2a: color = 2'b00;
		14'h0c2b: color = 2'b00;
		14'h0c2c: color = 2'b00;
		14'h0c2d: color = 2'b00;
		14'h0c2e: color = 2'b01;
		14'h0c2f: color = 2'b00;
		14'h0c30: color = 2'b00;
		14'h0c31: color = 2'b00;
		14'h0c32: color = 2'b00;
		14'h0c33: color = 2'b01;
		14'h0c34: color = 2'b00;
		14'h0c35: color = 2'b01;
		14'h0c36: color = 2'b00;
		14'h0c37: color = 2'b00;
		14'h0c38: color = 2'b00;
		14'h0c39: color = 2'b00;
		14'h0c3a: color = 2'b00;
		14'h0c3b: color = 2'b00;
		14'h0c3c: color = 2'b00;
		14'h0c3d: color = 2'b00;
		14'h0c3e: color = 2'b00;
		14'h0c3f: color = 2'b00;
		14'h0c40: color = 2'b00;
		14'h0c41: color = 2'b00;
		14'h0c42: color = 2'b00;
		14'h0c43: color = 2'b00;
		14'h0c44: color = 2'b00;
		14'h0c45: color = 2'b00;
		14'h0c46: color = 2'b00;
		14'h0c47: color = 2'b00;
		14'h0c48: color = 2'b00;
		14'h0c49: color = 2'b00;
		14'h0c4a: color = 2'b00;
		14'h0c4b: color = 2'b00;
		14'h0c4c: color = 2'b00;
		14'h0c4d: color = 2'b00;
		14'h0c4e: color = 2'b00;
		14'h0c4f: color = 2'b00;
		14'h0c50: color = 2'b00;
		14'h0c51: color = 2'b00;
		14'h0c52: color = 2'b00;
		14'h0c53: color = 2'b00;
		14'h0c54: color = 2'b00;
		14'h0c55: color = 2'b00;
		14'h0c56: color = 2'b00;
		14'h0c57: color = 2'b00;
		14'h0c58: color = 2'b00;
		14'h0c59: color = 2'b00;
		14'h0c5a: color = 2'b00;
		14'h0c5b: color = 2'b00;
		14'h0c5c: color = 2'b00;
		14'h0c5d: color = 2'b00;
		14'h0c5e: color = 2'b00;
		14'h0c5f: color = 2'b00;
		14'h0c60: color = 2'b00;
		14'h0c61: color = 2'b00;
		14'h0c62: color = 2'b00;
		14'h0c63: color = 2'b00;
		14'h0c64: color = 2'b00;
		14'h0c65: color = 2'b11;
		14'h0c66: color = 2'b11;
		14'h0c67: color = 2'b11;
		14'h0c68: color = 2'b11;
		14'h0c69: color = 2'b11;
		14'h0c6a: color = 2'b11;
		14'h0c6b: color = 2'b11;
		14'h0c6c: color = 2'b11;
		14'h0c6d: color = 2'b11;
		14'h0c6e: color = 2'b11;
		14'h0c6f: color = 2'b11;
		14'h0c70: color = 2'b11;
		14'h0c71: color = 2'b11;
		14'h0c72: color = 2'b11;
		14'h0c73: color = 2'b11;
		14'h0c74: color = 2'b11;
		14'h0c75: color = 2'b11;
		14'h0c76: color = 2'b11;
		14'h0c77: color = 2'b11;
		14'h0c78: color = 2'b11;
		14'h0c79: color = 2'b11;
		14'h0c7a: color = 2'b11;
		14'h0c7b: color = 2'b11;
		14'h0c7c: color = 2'b11;
		14'h0c7d: color = 2'b11;
		14'h0c7e: color = 2'b11;
		14'h0c7f: color = 2'b11;
		14'h0c80: color = 2'b11;
		14'h0c81: color = 2'b11;
		14'h0c82: color = 2'b11;
		14'h0c83: color = 2'b11;
		14'h0c84: color = 2'b11;
		14'h0c85: color = 2'b11;
		14'h0c86: color = 2'b11;
		14'h0c87: color = 2'b11;
		14'h0c88: color = 2'b11;
		14'h0c89: color = 2'b11;
		14'h0c8a: color = 2'b11;
		14'h0c8b: color = 2'b11;
		14'h0c8c: color = 2'b11;
		14'h0c8d: color = 2'b11;
		14'h0c8e: color = 2'b11;
		14'h0c8f: color = 2'b11;
		14'h0c90: color = 2'b11;
		14'h0c91: color = 2'b11;
		14'h0c92: color = 2'b11;
		14'h0c93: color = 2'b11;
		14'h0c94: color = 2'b11;
		14'h0c95: color = 2'b11;
		14'h0c96: color = 2'b11;
		14'h0c97: color = 2'b11;
		14'h0c98: color = 2'b11;
		14'h0c99: color = 2'b11;
		14'h0c9a: color = 2'b11;
		14'h0c9b: color = 2'b11;
		14'h0c9c: color = 2'b11;
		14'h0c9d: color = 2'b11;
		14'h0c9e: color = 2'b11;
		14'h0c9f: color = 2'b11;
		14'h0ca0: color = 2'b11;
		14'h0ca1: color = 2'b11;
		14'h0ca2: color = 2'b11;
		14'h0ca3: color = 2'b11;
		14'h0ca4: color = 2'b11;
		14'h0ca5: color = 2'b10;
		14'h0ca6: color = 2'b10;
		14'h0ca7: color = 2'b00;
		14'h0ca8: color = 2'b00;
		14'h0ca9: color = 2'b00;
		14'h0caa: color = 2'b00;
		14'h0cab: color = 2'b00;
		14'h0cac: color = 2'b00;
		14'h0cad: color = 2'b00;
		14'h0cae: color = 2'b00;
		14'h0caf: color = 2'b00;
		14'h0cb0: color = 2'b01;
		14'h0cb1: color = 2'b01;
		14'h0cb2: color = 2'b01;
		14'h0cb3: color = 2'b01;
		14'h0cb4: color = 2'b00;
		14'h0cb5: color = 2'b00;
		14'h0cb6: color = 2'b00;
		14'h0cb7: color = 2'b00;
		14'h0cb8: color = 2'b00;
		14'h0cb9: color = 2'b00;
		14'h0cba: color = 2'b00;
		14'h0cbb: color = 2'b00;
		14'h0cbc: color = 2'b00;
		14'h0cbd: color = 2'b00;
		14'h0cbe: color = 2'b00;
		14'h0cbf: color = 2'b00;
		14'h0cc0: color = 2'b00;
		14'h0cc1: color = 2'b00;
		14'h0cc2: color = 2'b00;
		14'h0cc3: color = 2'b00;
		14'h0cc4: color = 2'b00;
		14'h0cc5: color = 2'b00;
		14'h0cc6: color = 2'b00;
		14'h0cc7: color = 2'b00;
		14'h0cc8: color = 2'b00;
		14'h0cc9: color = 2'b00;
		14'h0cca: color = 2'b00;
		14'h0ccb: color = 2'b00;
		14'h0ccc: color = 2'b00;
		14'h0ccd: color = 2'b00;
		14'h0cce: color = 2'b00;
		14'h0ccf: color = 2'b00;
		14'h0cd0: color = 2'b00;
		14'h0cd1: color = 2'b00;
		14'h0cd2: color = 2'b00;
		14'h0cd3: color = 2'b00;
		14'h0cd4: color = 2'b00;
		14'h0cd5: color = 2'b00;
		14'h0cd6: color = 2'b00;
		14'h0cd7: color = 2'b00;
		14'h0cd8: color = 2'b00;
		14'h0cd9: color = 2'b00;
		14'h0cda: color = 2'b00;
		14'h0cdb: color = 2'b00;
		14'h0cdc: color = 2'b00;
		14'h0cdd: color = 2'b00;
		14'h0cde: color = 2'b00;
		14'h0cdf: color = 2'b00;
		14'h0ce0: color = 2'b00;
		14'h0ce1: color = 2'b00;
		14'h0ce2: color = 2'b00;
		14'h0ce3: color = 2'b00;
		14'h0ce4: color = 2'b00;
		14'h0ce5: color = 2'b01;
		14'h0ce6: color = 2'b11;
		14'h0ce7: color = 2'b11;
		14'h0ce8: color = 2'b11;
		14'h0ce9: color = 2'b11;
		14'h0cea: color = 2'b11;
		14'h0ceb: color = 2'b11;
		14'h0cec: color = 2'b11;
		14'h0ced: color = 2'b11;
		14'h0cee: color = 2'b11;
		14'h0cef: color = 2'b11;
		14'h0cf0: color = 2'b11;
		14'h0cf1: color = 2'b11;
		14'h0cf2: color = 2'b11;
		14'h0cf3: color = 2'b11;
		14'h0cf4: color = 2'b11;
		14'h0cf5: color = 2'b11;
		14'h0cf6: color = 2'b11;
		14'h0cf7: color = 2'b11;
		14'h0cf8: color = 2'b11;
		14'h0cf9: color = 2'b11;
		14'h0cfa: color = 2'b11;
		14'h0cfb: color = 2'b11;
		14'h0cfc: color = 2'b11;
		14'h0cfd: color = 2'b11;
		14'h0cfe: color = 2'b11;
		14'h0cff: color = 2'b11;
		14'h0d00: color = 2'b11;
		14'h0d01: color = 2'b11;
		14'h0d02: color = 2'b11;
		14'h0d03: color = 2'b11;
		14'h0d04: color = 2'b11;
		14'h0d05: color = 2'b11;
		14'h0d06: color = 2'b11;
		14'h0d07: color = 2'b11;
		14'h0d08: color = 2'b11;
		14'h0d09: color = 2'b11;
		14'h0d0a: color = 2'b11;
		14'h0d0b: color = 2'b11;
		14'h0d0c: color = 2'b11;
		14'h0d0d: color = 2'b11;
		14'h0d0e: color = 2'b11;
		14'h0d0f: color = 2'b11;
		14'h0d10: color = 2'b11;
		14'h0d11: color = 2'b11;
		14'h0d12: color = 2'b11;
		14'h0d13: color = 2'b11;
		14'h0d14: color = 2'b11;
		14'h0d15: color = 2'b11;
		14'h0d16: color = 2'b11;
		14'h0d17: color = 2'b11;
		14'h0d18: color = 2'b11;
		14'h0d19: color = 2'b11;
		14'h0d1a: color = 2'b11;
		14'h0d1b: color = 2'b11;
		14'h0d1c: color = 2'b11;
		14'h0d1d: color = 2'b11;
		14'h0d1e: color = 2'b11;
		14'h0d1f: color = 2'b11;
		14'h0d20: color = 2'b11;
		14'h0d21: color = 2'b11;
		14'h0d22: color = 2'b11;
		14'h0d23: color = 2'b11;
		14'h0d24: color = 2'b11;
		14'h0d25: color = 2'b00;
		14'h0d26: color = 2'b00;
		14'h0d27: color = 2'b00;
		14'h0d28: color = 2'b00;
		14'h0d29: color = 2'b00;
		14'h0d2a: color = 2'b00;
		14'h0d2b: color = 2'b00;
		14'h0d2c: color = 2'b00;
		14'h0d2d: color = 2'b01;
		14'h0d2e: color = 2'b01;
		14'h0d2f: color = 2'b01;
		14'h0d30: color = 2'b00;
		14'h0d31: color = 2'b00;
		14'h0d32: color = 2'b01;
		14'h0d33: color = 2'b00;
		14'h0d34: color = 2'b00;
		14'h0d35: color = 2'b00;
		14'h0d36: color = 2'b00;
		14'h0d37: color = 2'b00;
		14'h0d38: color = 2'b00;
		14'h0d39: color = 2'b00;
		14'h0d3a: color = 2'b00;
		14'h0d3b: color = 2'b00;
		14'h0d3c: color = 2'b00;
		14'h0d3d: color = 2'b00;
		14'h0d3e: color = 2'b00;
		14'h0d3f: color = 2'b00;
		14'h0d40: color = 2'b00;
		14'h0d41: color = 2'b00;
		14'h0d42: color = 2'b00;
		14'h0d43: color = 2'b00;
		14'h0d44: color = 2'b00;
		14'h0d45: color = 2'b00;
		14'h0d46: color = 2'b00;
		14'h0d47: color = 2'b00;
		14'h0d48: color = 2'b00;
		14'h0d49: color = 2'b00;
		14'h0d4a: color = 2'b00;
		14'h0d4b: color = 2'b00;
		14'h0d4c: color = 2'b00;
		14'h0d4d: color = 2'b00;
		14'h0d4e: color = 2'b00;
		14'h0d4f: color = 2'b00;
		14'h0d50: color = 2'b00;
		14'h0d51: color = 2'b00;
		14'h0d52: color = 2'b00;
		14'h0d53: color = 2'b00;
		14'h0d54: color = 2'b00;
		14'h0d55: color = 2'b00;
		14'h0d56: color = 2'b00;
		14'h0d57: color = 2'b00;
		14'h0d58: color = 2'b00;
		14'h0d59: color = 2'b00;
		14'h0d5a: color = 2'b00;
		14'h0d5b: color = 2'b00;
		14'h0d5c: color = 2'b00;
		14'h0d5d: color = 2'b00;
		14'h0d5e: color = 2'b00;
		14'h0d5f: color = 2'b00;
		14'h0d60: color = 2'b00;
		14'h0d61: color = 2'b00;
		14'h0d62: color = 2'b00;
		14'h0d63: color = 2'b00;
		14'h0d64: color = 2'b00;
		14'h0d65: color = 2'b00;
		14'h0d66: color = 2'b11;
		14'h0d67: color = 2'b11;
		14'h0d68: color = 2'b11;
		14'h0d69: color = 2'b11;
		14'h0d6a: color = 2'b11;
		14'h0d6b: color = 2'b11;
		14'h0d6c: color = 2'b11;
		14'h0d6d: color = 2'b11;
		14'h0d6e: color = 2'b11;
		14'h0d6f: color = 2'b11;
		14'h0d70: color = 2'b11;
		14'h0d71: color = 2'b11;
		14'h0d72: color = 2'b11;
		14'h0d73: color = 2'b11;
		14'h0d74: color = 2'b11;
		14'h0d75: color = 2'b11;
		14'h0d76: color = 2'b11;
		14'h0d77: color = 2'b11;
		14'h0d78: color = 2'b11;
		14'h0d79: color = 2'b11;
		14'h0d7a: color = 2'b11;
		14'h0d7b: color = 2'b11;
		14'h0d7c: color = 2'b11;
		14'h0d7d: color = 2'b11;
		14'h0d7e: color = 2'b11;
		14'h0d7f: color = 2'b11;
		14'h0d80: color = 2'b11;
		14'h0d81: color = 2'b11;
		14'h0d82: color = 2'b11;
		14'h0d83: color = 2'b11;
		14'h0d84: color = 2'b11;
		14'h0d85: color = 2'b11;
		14'h0d86: color = 2'b11;
		14'h0d87: color = 2'b11;
		14'h0d88: color = 2'b11;
		14'h0d89: color = 2'b11;
		14'h0d8a: color = 2'b11;
		14'h0d8b: color = 2'b11;
		14'h0d8c: color = 2'b11;
		14'h0d8d: color = 2'b11;
		14'h0d8e: color = 2'b11;
		14'h0d8f: color = 2'b11;
		14'h0d90: color = 2'b11;
		14'h0d91: color = 2'b11;
		14'h0d92: color = 2'b11;
		14'h0d93: color = 2'b11;
		14'h0d94: color = 2'b11;
		14'h0d95: color = 2'b11;
		14'h0d96: color = 2'b11;
		14'h0d97: color = 2'b11;
		14'h0d98: color = 2'b11;
		14'h0d99: color = 2'b11;
		14'h0d9a: color = 2'b11;
		14'h0d9b: color = 2'b11;
		14'h0d9c: color = 2'b11;
		14'h0d9d: color = 2'b11;
		14'h0d9e: color = 2'b11;
		14'h0d9f: color = 2'b11;
		14'h0da0: color = 2'b11;
		14'h0da1: color = 2'b11;
		14'h0da2: color = 2'b11;
		14'h0da3: color = 2'b11;
		14'h0da4: color = 2'b01;
		14'h0da5: color = 2'b00;
		14'h0da6: color = 2'b00;
		14'h0da7: color = 2'b00;
		14'h0da8: color = 2'b00;
		14'h0da9: color = 2'b00;
		14'h0daa: color = 2'b00;
		14'h0dab: color = 2'b01;
		14'h0dac: color = 2'b01;
		14'h0dad: color = 2'b00;
		14'h0dae: color = 2'b01;
		14'h0daf: color = 2'b00;
		14'h0db0: color = 2'b00;
		14'h0db1: color = 2'b01;
		14'h0db2: color = 2'b01;
		14'h0db3: color = 2'b00;
		14'h0db4: color = 2'b00;
		14'h0db5: color = 2'b00;
		14'h0db6: color = 2'b00;
		14'h0db7: color = 2'b00;
		14'h0db8: color = 2'b00;
		14'h0db9: color = 2'b00;
		14'h0dba: color = 2'b00;
		14'h0dbb: color = 2'b00;
		14'h0dbc: color = 2'b00;
		14'h0dbd: color = 2'b00;
		14'h0dbe: color = 2'b00;
		14'h0dbf: color = 2'b00;
		14'h0dc0: color = 2'b00;
		14'h0dc1: color = 2'b00;
		14'h0dc2: color = 2'b00;
		14'h0dc3: color = 2'b00;
		14'h0dc4: color = 2'b00;
		14'h0dc5: color = 2'b00;
		14'h0dc6: color = 2'b00;
		14'h0dc7: color = 2'b00;
		14'h0dc8: color = 2'b00;
		14'h0dc9: color = 2'b00;
		14'h0dca: color = 2'b00;
		14'h0dcb: color = 2'b00;
		14'h0dcc: color = 2'b00;
		14'h0dcd: color = 2'b00;
		14'h0dce: color = 2'b00;
		14'h0dcf: color = 2'b00;
		14'h0dd0: color = 2'b00;
		14'h0dd1: color = 2'b00;
		14'h0dd2: color = 2'b00;
		14'h0dd3: color = 2'b00;
		14'h0dd4: color = 2'b00;
		14'h0dd5: color = 2'b00;
		14'h0dd6: color = 2'b00;
		14'h0dd7: color = 2'b00;
		14'h0dd8: color = 2'b00;
		14'h0dd9: color = 2'b00;
		14'h0dda: color = 2'b00;
		14'h0ddb: color = 2'b00;
		14'h0ddc: color = 2'b00;
		14'h0ddd: color = 2'b00;
		14'h0dde: color = 2'b00;
		14'h0ddf: color = 2'b00;
		14'h0de0: color = 2'b00;
		14'h0de1: color = 2'b00;
		14'h0de2: color = 2'b00;
		14'h0de3: color = 2'b00;
		14'h0de4: color = 2'b00;
		14'h0de5: color = 2'b00;
		14'h0de6: color = 2'b11;
		14'h0de7: color = 2'b11;
		14'h0de8: color = 2'b11;
		14'h0de9: color = 2'b11;
		14'h0dea: color = 2'b11;
		14'h0deb: color = 2'b11;
		14'h0dec: color = 2'b11;
		14'h0ded: color = 2'b11;
		14'h0dee: color = 2'b11;
		14'h0def: color = 2'b11;
		14'h0df0: color = 2'b11;
		14'h0df1: color = 2'b11;
		14'h0df2: color = 2'b11;
		14'h0df3: color = 2'b11;
		14'h0df4: color = 2'b11;
		14'h0df5: color = 2'b11;
		14'h0df6: color = 2'b11;
		14'h0df7: color = 2'b11;
		14'h0df8: color = 2'b11;
		14'h0df9: color = 2'b11;
		14'h0dfa: color = 2'b11;
		14'h0dfb: color = 2'b11;
		14'h0dfc: color = 2'b11;
		14'h0dfd: color = 2'b11;
		14'h0dfe: color = 2'b11;
		14'h0dff: color = 2'b11;
		14'h0e00: color = 2'b11;
		14'h0e01: color = 2'b11;
		14'h0e02: color = 2'b11;
		14'h0e03: color = 2'b11;
		14'h0e04: color = 2'b11;
		14'h0e05: color = 2'b11;
		14'h0e06: color = 2'b11;
		14'h0e07: color = 2'b11;
		14'h0e08: color = 2'b11;
		14'h0e09: color = 2'b11;
		14'h0e0a: color = 2'b11;
		14'h0e0b: color = 2'b11;
		14'h0e0c: color = 2'b11;
		14'h0e0d: color = 2'b11;
		14'h0e0e: color = 2'b11;
		14'h0e0f: color = 2'b11;
		14'h0e10: color = 2'b11;
		14'h0e11: color = 2'b11;
		14'h0e12: color = 2'b11;
		14'h0e13: color = 2'b11;
		14'h0e14: color = 2'b11;
		14'h0e15: color = 2'b11;
		14'h0e16: color = 2'b11;
		14'h0e17: color = 2'b11;
		14'h0e18: color = 2'b11;
		14'h0e19: color = 2'b11;
		14'h0e1a: color = 2'b11;
		14'h0e1b: color = 2'b11;
		14'h0e1c: color = 2'b11;
		14'h0e1d: color = 2'b11;
		14'h0e1e: color = 2'b11;
		14'h0e1f: color = 2'b11;
		14'h0e20: color = 2'b11;
		14'h0e21: color = 2'b11;
		14'h0e22: color = 2'b11;
		14'h0e23: color = 2'b11;
		14'h0e24: color = 2'b00;
		14'h0e25: color = 2'b00;
		14'h0e26: color = 2'b00;
		14'h0e27: color = 2'b00;
		14'h0e28: color = 2'b00;
		14'h0e29: color = 2'b00;
		14'h0e2a: color = 2'b01;
		14'h0e2b: color = 2'b00;
		14'h0e2c: color = 2'b01;
		14'h0e2d: color = 2'b00;
		14'h0e2e: color = 2'b01;
		14'h0e2f: color = 2'b01;
		14'h0e30: color = 2'b00;
		14'h0e31: color = 2'b00;
		14'h0e32: color = 2'b01;
		14'h0e33: color = 2'b01;
		14'h0e34: color = 2'b00;
		14'h0e35: color = 2'b00;
		14'h0e36: color = 2'b00;
		14'h0e37: color = 2'b00;
		14'h0e38: color = 2'b00;
		14'h0e39: color = 2'b00;
		14'h0e3a: color = 2'b00;
		14'h0e3b: color = 2'b01;
		14'h0e3c: color = 2'b00;
		14'h0e3d: color = 2'b00;
		14'h0e3e: color = 2'b00;
		14'h0e3f: color = 2'b00;
		14'h0e40: color = 2'b00;
		14'h0e41: color = 2'b00;
		14'h0e42: color = 2'b00;
		14'h0e43: color = 2'b00;
		14'h0e44: color = 2'b00;
		14'h0e45: color = 2'b00;
		14'h0e46: color = 2'b00;
		14'h0e47: color = 2'b00;
		14'h0e48: color = 2'b00;
		14'h0e49: color = 2'b00;
		14'h0e4a: color = 2'b00;
		14'h0e4b: color = 2'b00;
		14'h0e4c: color = 2'b00;
		14'h0e4d: color = 2'b00;
		14'h0e4e: color = 2'b00;
		14'h0e4f: color = 2'b00;
		14'h0e50: color = 2'b00;
		14'h0e51: color = 2'b00;
		14'h0e52: color = 2'b00;
		14'h0e53: color = 2'b00;
		14'h0e54: color = 2'b00;
		14'h0e55: color = 2'b00;
		14'h0e56: color = 2'b00;
		14'h0e57: color = 2'b00;
		14'h0e58: color = 2'b00;
		14'h0e59: color = 2'b00;
		14'h0e5a: color = 2'b00;
		14'h0e5b: color = 2'b00;
		14'h0e5c: color = 2'b00;
		14'h0e5d: color = 2'b00;
		14'h0e5e: color = 2'b00;
		14'h0e5f: color = 2'b00;
		14'h0e60: color = 2'b00;
		14'h0e61: color = 2'b00;
		14'h0e62: color = 2'b00;
		14'h0e63: color = 2'b00;
		14'h0e64: color = 2'b00;
		14'h0e65: color = 2'b00;
		14'h0e66: color = 2'b01;
		14'h0e67: color = 2'b11;
		14'h0e68: color = 2'b11;
		14'h0e69: color = 2'b11;
		14'h0e6a: color = 2'b11;
		14'h0e6b: color = 2'b11;
		14'h0e6c: color = 2'b11;
		14'h0e6d: color = 2'b11;
		14'h0e6e: color = 2'b11;
		14'h0e6f: color = 2'b11;
		14'h0e70: color = 2'b11;
		14'h0e71: color = 2'b11;
		14'h0e72: color = 2'b11;
		14'h0e73: color = 2'b11;
		14'h0e74: color = 2'b11;
		14'h0e75: color = 2'b11;
		14'h0e76: color = 2'b11;
		14'h0e77: color = 2'b11;
		14'h0e78: color = 2'b11;
		14'h0e79: color = 2'b11;
		14'h0e7a: color = 2'b11;
		14'h0e7b: color = 2'b11;
		14'h0e7c: color = 2'b11;
		14'h0e7d: color = 2'b11;
		14'h0e7e: color = 2'b11;
		14'h0e7f: color = 2'b11;
		14'h0e80: color = 2'b11;
		14'h0e81: color = 2'b11;
		14'h0e82: color = 2'b11;
		14'h0e83: color = 2'b11;
		14'h0e84: color = 2'b11;
		14'h0e85: color = 2'b11;
		14'h0e86: color = 2'b11;
		14'h0e87: color = 2'b11;
		14'h0e88: color = 2'b11;
		14'h0e89: color = 2'b11;
		14'h0e8a: color = 2'b11;
		14'h0e8b: color = 2'b11;
		14'h0e8c: color = 2'b11;
		14'h0e8d: color = 2'b11;
		14'h0e8e: color = 2'b11;
		14'h0e8f: color = 2'b11;
		14'h0e90: color = 2'b11;
		14'h0e91: color = 2'b11;
		14'h0e92: color = 2'b11;
		14'h0e93: color = 2'b11;
		14'h0e94: color = 2'b11;
		14'h0e95: color = 2'b11;
		14'h0e96: color = 2'b11;
		14'h0e97: color = 2'b11;
		14'h0e98: color = 2'b11;
		14'h0e99: color = 2'b11;
		14'h0e9a: color = 2'b11;
		14'h0e9b: color = 2'b11;
		14'h0e9c: color = 2'b11;
		14'h0e9d: color = 2'b11;
		14'h0e9e: color = 2'b11;
		14'h0e9f: color = 2'b11;
		14'h0ea0: color = 2'b11;
		14'h0ea1: color = 2'b11;
		14'h0ea2: color = 2'b11;
		14'h0ea3: color = 2'b11;
		14'h0ea4: color = 2'b00;
		14'h0ea5: color = 2'b01;
		14'h0ea6: color = 2'b00;
		14'h0ea7: color = 2'b01;
		14'h0ea8: color = 2'b01;
		14'h0ea9: color = 2'b00;
		14'h0eaa: color = 2'b01;
		14'h0eab: color = 2'b00;
		14'h0eac: color = 2'b00;
		14'h0ead: color = 2'b01;
		14'h0eae: color = 2'b00;
		14'h0eaf: color = 2'b01;
		14'h0eb0: color = 2'b00;
		14'h0eb1: color = 2'b01;
		14'h0eb2: color = 2'b00;
		14'h0eb3: color = 2'b01;
		14'h0eb4: color = 2'b00;
		14'h0eb5: color = 2'b00;
		14'h0eb6: color = 2'b00;
		14'h0eb7: color = 2'b00;
		14'h0eb8: color = 2'b00;
		14'h0eb9: color = 2'b00;
		14'h0eba: color = 2'b00;
		14'h0ebb: color = 2'b00;
		14'h0ebc: color = 2'b00;
		14'h0ebd: color = 2'b01;
		14'h0ebe: color = 2'b00;
		14'h0ebf: color = 2'b00;
		14'h0ec0: color = 2'b00;
		14'h0ec1: color = 2'b00;
		14'h0ec2: color = 2'b00;
		14'h0ec3: color = 2'b00;
		14'h0ec4: color = 2'b00;
		14'h0ec5: color = 2'b00;
		14'h0ec6: color = 2'b00;
		14'h0ec7: color = 2'b00;
		14'h0ec8: color = 2'b00;
		14'h0ec9: color = 2'b00;
		14'h0eca: color = 2'b00;
		14'h0ecb: color = 2'b00;
		14'h0ecc: color = 2'b00;
		14'h0ecd: color = 2'b00;
		14'h0ece: color = 2'b00;
		14'h0ecf: color = 2'b00;
		14'h0ed0: color = 2'b00;
		14'h0ed1: color = 2'b00;
		14'h0ed2: color = 2'b00;
		14'h0ed3: color = 2'b00;
		14'h0ed4: color = 2'b00;
		14'h0ed5: color = 2'b00;
		14'h0ed6: color = 2'b00;
		14'h0ed7: color = 2'b00;
		14'h0ed8: color = 2'b00;
		14'h0ed9: color = 2'b00;
		14'h0eda: color = 2'b00;
		14'h0edb: color = 2'b00;
		14'h0edc: color = 2'b00;
		14'h0edd: color = 2'b00;
		14'h0ede: color = 2'b00;
		14'h0edf: color = 2'b00;
		14'h0ee0: color = 2'b00;
		14'h0ee1: color = 2'b00;
		14'h0ee2: color = 2'b00;
		14'h0ee3: color = 2'b00;
		14'h0ee4: color = 2'b00;
		14'h0ee5: color = 2'b00;
		14'h0ee6: color = 2'b00;
		14'h0ee7: color = 2'b11;
		14'h0ee8: color = 2'b11;
		14'h0ee9: color = 2'b11;
		14'h0eea: color = 2'b11;
		14'h0eeb: color = 2'b11;
		14'h0eec: color = 2'b11;
		14'h0eed: color = 2'b11;
		14'h0eee: color = 2'b11;
		14'h0eef: color = 2'b11;
		14'h0ef0: color = 2'b11;
		14'h0ef1: color = 2'b11;
		14'h0ef2: color = 2'b11;
		14'h0ef3: color = 2'b11;
		14'h0ef4: color = 2'b11;
		14'h0ef5: color = 2'b11;
		14'h0ef6: color = 2'b11;
		14'h0ef7: color = 2'b11;
		14'h0ef8: color = 2'b11;
		14'h0ef9: color = 2'b11;
		14'h0efa: color = 2'b11;
		14'h0efb: color = 2'b11;
		14'h0efc: color = 2'b11;
		14'h0efd: color = 2'b11;
		14'h0efe: color = 2'b11;
		14'h0eff: color = 2'b11;
		14'h0f00: color = 2'b11;
		14'h0f01: color = 2'b11;
		14'h0f02: color = 2'b11;
		14'h0f03: color = 2'b11;
		14'h0f04: color = 2'b11;
		14'h0f05: color = 2'b11;
		14'h0f06: color = 2'b11;
		14'h0f07: color = 2'b11;
		14'h0f08: color = 2'b11;
		14'h0f09: color = 2'b11;
		14'h0f0a: color = 2'b11;
		14'h0f0b: color = 2'b11;
		14'h0f0c: color = 2'b11;
		14'h0f0d: color = 2'b11;
		14'h0f0e: color = 2'b11;
		14'h0f0f: color = 2'b11;
		14'h0f10: color = 2'b11;
		14'h0f11: color = 2'b11;
		14'h0f12: color = 2'b11;
		14'h0f13: color = 2'b11;
		14'h0f14: color = 2'b11;
		14'h0f15: color = 2'b11;
		14'h0f16: color = 2'b11;
		14'h0f17: color = 2'b11;
		14'h0f18: color = 2'b11;
		14'h0f19: color = 2'b11;
		14'h0f1a: color = 2'b11;
		14'h0f1b: color = 2'b11;
		14'h0f1c: color = 2'b11;
		14'h0f1d: color = 2'b11;
		14'h0f1e: color = 2'b11;
		14'h0f1f: color = 2'b11;
		14'h0f20: color = 2'b11;
		14'h0f21: color = 2'b11;
		14'h0f22: color = 2'b11;
		14'h0f23: color = 2'b10;
		14'h0f24: color = 2'b00;
		14'h0f25: color = 2'b00;
		14'h0f26: color = 2'b00;
		14'h0f27: color = 2'b00;
		14'h0f28: color = 2'b00;
		14'h0f29: color = 2'b00;
		14'h0f2a: color = 2'b01;
		14'h0f2b: color = 2'b01;
		14'h0f2c: color = 2'b00;
		14'h0f2d: color = 2'b00;
		14'h0f2e: color = 2'b01;
		14'h0f2f: color = 2'b00;
		14'h0f30: color = 2'b00;
		14'h0f31: color = 2'b01;
		14'h0f32: color = 2'b00;
		14'h0f33: color = 2'b00;
		14'h0f34: color = 2'b00;
		14'h0f35: color = 2'b00;
		14'h0f36: color = 2'b00;
		14'h0f37: color = 2'b00;
		14'h0f38: color = 2'b00;
		14'h0f39: color = 2'b00;
		14'h0f3a: color = 2'b00;
		14'h0f3b: color = 2'b01;
		14'h0f3c: color = 2'b00;
		14'h0f3d: color = 2'b00;
		14'h0f3e: color = 2'b01;
		14'h0f3f: color = 2'b00;
		14'h0f40: color = 2'b00;
		14'h0f41: color = 2'b00;
		14'h0f42: color = 2'b00;
		14'h0f43: color = 2'b00;
		14'h0f44: color = 2'b00;
		14'h0f45: color = 2'b00;
		14'h0f46: color = 2'b00;
		14'h0f47: color = 2'b00;
		14'h0f48: color = 2'b00;
		14'h0f49: color = 2'b00;
		14'h0f4a: color = 2'b00;
		14'h0f4b: color = 2'b00;
		14'h0f4c: color = 2'b00;
		14'h0f4d: color = 2'b00;
		14'h0f4e: color = 2'b00;
		14'h0f4f: color = 2'b00;
		14'h0f50: color = 2'b00;
		14'h0f51: color = 2'b00;
		14'h0f52: color = 2'b00;
		14'h0f53: color = 2'b00;
		14'h0f54: color = 2'b00;
		14'h0f55: color = 2'b00;
		14'h0f56: color = 2'b00;
		14'h0f57: color = 2'b00;
		14'h0f58: color = 2'b00;
		14'h0f59: color = 2'b00;
		14'h0f5a: color = 2'b00;
		14'h0f5b: color = 2'b01;
		14'h0f5c: color = 2'b01;
		14'h0f5d: color = 2'b00;
		14'h0f5e: color = 2'b00;
		14'h0f5f: color = 2'b00;
		14'h0f60: color = 2'b00;
		14'h0f61: color = 2'b00;
		14'h0f62: color = 2'b00;
		14'h0f63: color = 2'b00;
		14'h0f64: color = 2'b00;
		14'h0f65: color = 2'b00;
		14'h0f66: color = 2'b00;
		14'h0f67: color = 2'b11;
		14'h0f68: color = 2'b11;
		14'h0f69: color = 2'b11;
		14'h0f6a: color = 2'b11;
		14'h0f6b: color = 2'b11;
		14'h0f6c: color = 2'b11;
		14'h0f6d: color = 2'b11;
		14'h0f6e: color = 2'b11;
		14'h0f6f: color = 2'b11;
		14'h0f70: color = 2'b11;
		14'h0f71: color = 2'b11;
		14'h0f72: color = 2'b11;
		14'h0f73: color = 2'b11;
		14'h0f74: color = 2'b11;
		14'h0f75: color = 2'b11;
		14'h0f76: color = 2'b11;
		14'h0f77: color = 2'b11;
		14'h0f78: color = 2'b11;
		14'h0f79: color = 2'b11;
		14'h0f7a: color = 2'b11;
		14'h0f7b: color = 2'b11;
		14'h0f7c: color = 2'b11;
		14'h0f7d: color = 2'b11;
		14'h0f7e: color = 2'b11;
		14'h0f7f: color = 2'b11;
		14'h0f80: color = 2'b11;
		14'h0f81: color = 2'b11;
		14'h0f82: color = 2'b11;
		14'h0f83: color = 2'b11;
		14'h0f84: color = 2'b11;
		14'h0f85: color = 2'b11;
		14'h0f86: color = 2'b11;
		14'h0f87: color = 2'b11;
		14'h0f88: color = 2'b11;
		14'h0f89: color = 2'b11;
		14'h0f8a: color = 2'b11;
		14'h0f8b: color = 2'b11;
		14'h0f8c: color = 2'b11;
		14'h0f8d: color = 2'b11;
		14'h0f8e: color = 2'b11;
		14'h0f8f: color = 2'b11;
		14'h0f90: color = 2'b11;
		14'h0f91: color = 2'b11;
		14'h0f92: color = 2'b11;
		14'h0f93: color = 2'b11;
		14'h0f94: color = 2'b11;
		14'h0f95: color = 2'b11;
		14'h0f96: color = 2'b11;
		14'h0f97: color = 2'b11;
		14'h0f98: color = 2'b11;
		14'h0f99: color = 2'b11;
		14'h0f9a: color = 2'b11;
		14'h0f9b: color = 2'b11;
		14'h0f9c: color = 2'b11;
		14'h0f9d: color = 2'b11;
		14'h0f9e: color = 2'b11;
		14'h0f9f: color = 2'b11;
		14'h0fa0: color = 2'b11;
		14'h0fa1: color = 2'b11;
		14'h0fa2: color = 2'b11;
		14'h0fa3: color = 2'b01;
		14'h0fa4: color = 2'b00;
		14'h0fa5: color = 2'b00;
		14'h0fa6: color = 2'b00;
		14'h0fa7: color = 2'b00;
		14'h0fa8: color = 2'b00;
		14'h0fa9: color = 2'b00;
		14'h0faa: color = 2'b01;
		14'h0fab: color = 2'b00;
		14'h0fac: color = 2'b01;
		14'h0fad: color = 2'b00;
		14'h0fae: color = 2'b00;
		14'h0faf: color = 2'b01;
		14'h0fb0: color = 2'b01;
		14'h0fb1: color = 2'b00;
		14'h0fb2: color = 2'b01;
		14'h0fb3: color = 2'b00;
		14'h0fb4: color = 2'b00;
		14'h0fb5: color = 2'b00;
		14'h0fb6: color = 2'b00;
		14'h0fb7: color = 2'b00;
		14'h0fb8: color = 2'b00;
		14'h0fb9: color = 2'b01;
		14'h0fba: color = 2'b00;
		14'h0fbb: color = 2'b00;
		14'h0fbc: color = 2'b00;
		14'h0fbd: color = 2'b01;
		14'h0fbe: color = 2'b00;
		14'h0fbf: color = 2'b01;
		14'h0fc0: color = 2'b00;
		14'h0fc1: color = 2'b00;
		14'h0fc2: color = 2'b00;
		14'h0fc3: color = 2'b00;
		14'h0fc4: color = 2'b00;
		14'h0fc5: color = 2'b00;
		14'h0fc6: color = 2'b00;
		14'h0fc7: color = 2'b00;
		14'h0fc8: color = 2'b00;
		14'h0fc9: color = 2'b00;
		14'h0fca: color = 2'b00;
		14'h0fcb: color = 2'b00;
		14'h0fcc: color = 2'b00;
		14'h0fcd: color = 2'b00;
		14'h0fce: color = 2'b00;
		14'h0fcf: color = 2'b00;
		14'h0fd0: color = 2'b00;
		14'h0fd1: color = 2'b00;
		14'h0fd2: color = 2'b00;
		14'h0fd3: color = 2'b00;
		14'h0fd4: color = 2'b00;
		14'h0fd5: color = 2'b00;
		14'h0fd6: color = 2'b00;
		14'h0fd7: color = 2'b00;
		14'h0fd8: color = 2'b00;
		14'h0fd9: color = 2'b01;
		14'h0fda: color = 2'b01;
		14'h0fdb: color = 2'b01;
		14'h0fdc: color = 2'b01;
		14'h0fdd: color = 2'b01;
		14'h0fde: color = 2'b00;
		14'h0fdf: color = 2'b00;
		14'h0fe0: color = 2'b00;
		14'h0fe1: color = 2'b00;
		14'h0fe2: color = 2'b00;
		14'h0fe3: color = 2'b00;
		14'h0fe4: color = 2'b00;
		14'h0fe5: color = 2'b00;
		14'h0fe6: color = 2'b00;
		14'h0fe7: color = 2'b11;
		14'h0fe8: color = 2'b11;
		14'h0fe9: color = 2'b11;
		14'h0fea: color = 2'b11;
		14'h0feb: color = 2'b11;
		14'h0fec: color = 2'b11;
		14'h0fed: color = 2'b11;
		14'h0fee: color = 2'b11;
		14'h0fef: color = 2'b11;
		14'h0ff0: color = 2'b11;
		14'h0ff1: color = 2'b11;
		14'h0ff2: color = 2'b11;
		14'h0ff3: color = 2'b11;
		14'h0ff4: color = 2'b11;
		14'h0ff5: color = 2'b11;
		14'h0ff6: color = 2'b11;
		14'h0ff7: color = 2'b11;
		14'h0ff8: color = 2'b11;
		14'h0ff9: color = 2'b11;
		14'h0ffa: color = 2'b11;
		14'h0ffb: color = 2'b11;
		14'h0ffc: color = 2'b11;
		14'h0ffd: color = 2'b11;
		14'h0ffe: color = 2'b11;
		14'h0fff: color = 2'b11;
		14'h1000: color = 2'b11;
		14'h1001: color = 2'b11;
		14'h1002: color = 2'b11;
		14'h1003: color = 2'b11;
		14'h1004: color = 2'b11;
		14'h1005: color = 2'b11;
		14'h1006: color = 2'b11;
		14'h1007: color = 2'b11;
		14'h1008: color = 2'b11;
		14'h1009: color = 2'b11;
		14'h100a: color = 2'b11;
		14'h100b: color = 2'b11;
		14'h100c: color = 2'b11;
		14'h100d: color = 2'b11;
		14'h100e: color = 2'b11;
		14'h100f: color = 2'b11;
		14'h1010: color = 2'b11;
		14'h1011: color = 2'b11;
		14'h1012: color = 2'b11;
		14'h1013: color = 2'b11;
		14'h1014: color = 2'b11;
		14'h1015: color = 2'b11;
		14'h1016: color = 2'b11;
		14'h1017: color = 2'b11;
		14'h1018: color = 2'b11;
		14'h1019: color = 2'b11;
		14'h101a: color = 2'b11;
		14'h101b: color = 2'b11;
		14'h101c: color = 2'b11;
		14'h101d: color = 2'b11;
		14'h101e: color = 2'b11;
		14'h101f: color = 2'b11;
		14'h1020: color = 2'b11;
		14'h1021: color = 2'b11;
		14'h1022: color = 2'b11;
		14'h1023: color = 2'b01;
		14'h1024: color = 2'b00;
		14'h1025: color = 2'b00;
		14'h1026: color = 2'b00;
		14'h1027: color = 2'b00;
		14'h1028: color = 2'b00;
		14'h1029: color = 2'b01;
		14'h102a: color = 2'b00;
		14'h102b: color = 2'b01;
		14'h102c: color = 2'b01;
		14'h102d: color = 2'b01;
		14'h102e: color = 2'b00;
		14'h102f: color = 2'b00;
		14'h1030: color = 2'b00;
		14'h1031: color = 2'b00;
		14'h1032: color = 2'b00;
		14'h1033: color = 2'b00;
		14'h1034: color = 2'b00;
		14'h1035: color = 2'b00;
		14'h1036: color = 2'b00;
		14'h1037: color = 2'b00;
		14'h1038: color = 2'b00;
		14'h1039: color = 2'b00;
		14'h103a: color = 2'b00;
		14'h103b: color = 2'b00;
		14'h103c: color = 2'b00;
		14'h103d: color = 2'b00;
		14'h103e: color = 2'b00;
		14'h103f: color = 2'b01;
		14'h1040: color = 2'b00;
		14'h1041: color = 2'b00;
		14'h1042: color = 2'b00;
		14'h1043: color = 2'b00;
		14'h1044: color = 2'b00;
		14'h1045: color = 2'b00;
		14'h1046: color = 2'b00;
		14'h1047: color = 2'b00;
		14'h1048: color = 2'b00;
		14'h1049: color = 2'b00;
		14'h104a: color = 2'b00;
		14'h104b: color = 2'b00;
		14'h104c: color = 2'b00;
		14'h104d: color = 2'b00;
		14'h104e: color = 2'b00;
		14'h104f: color = 2'b00;
		14'h1050: color = 2'b00;
		14'h1051: color = 2'b00;
		14'h1052: color = 2'b00;
		14'h1053: color = 2'b00;
		14'h1054: color = 2'b00;
		14'h1055: color = 2'b01;
		14'h1056: color = 2'b01;
		14'h1057: color = 2'b01;
		14'h1058: color = 2'b01;
		14'h1059: color = 2'b01;
		14'h105a: color = 2'b01;
		14'h105b: color = 2'b01;
		14'h105c: color = 2'b01;
		14'h105d: color = 2'b01;
		14'h105e: color = 2'b01;
		14'h105f: color = 2'b00;
		14'h1060: color = 2'b00;
		14'h1061: color = 2'b00;
		14'h1062: color = 2'b00;
		14'h1063: color = 2'b00;
		14'h1064: color = 2'b00;
		14'h1065: color = 2'b00;
		14'h1066: color = 2'b00;
		14'h1067: color = 2'b10;
		14'h1068: color = 2'b10;
		14'h1069: color = 2'b11;
		14'h106a: color = 2'b11;
		14'h106b: color = 2'b11;
		14'h106c: color = 2'b11;
		14'h106d: color = 2'b11;
		14'h106e: color = 2'b11;
		14'h106f: color = 2'b11;
		14'h1070: color = 2'b11;
		14'h1071: color = 2'b11;
		14'h1072: color = 2'b11;
		14'h1073: color = 2'b11;
		14'h1074: color = 2'b11;
		14'h1075: color = 2'b11;
		14'h1076: color = 2'b11;
		14'h1077: color = 2'b11;
		14'h1078: color = 2'b11;
		14'h1079: color = 2'b11;
		14'h107a: color = 2'b11;
		14'h107b: color = 2'b11;
		14'h107c: color = 2'b11;
		14'h107d: color = 2'b11;
		14'h107e: color = 2'b11;
		14'h107f: color = 2'b11;
		14'h1080: color = 2'b11;
		14'h1081: color = 2'b11;
		14'h1082: color = 2'b11;
		14'h1083: color = 2'b11;
		14'h1084: color = 2'b11;
		14'h1085: color = 2'b11;
		14'h1086: color = 2'b11;
		14'h1087: color = 2'b11;
		14'h1088: color = 2'b11;
		14'h1089: color = 2'b11;
		14'h108a: color = 2'b11;
		14'h108b: color = 2'b11;
		14'h108c: color = 2'b11;
		14'h108d: color = 2'b11;
		14'h108e: color = 2'b11;
		14'h108f: color = 2'b11;
		14'h1090: color = 2'b11;
		14'h1091: color = 2'b11;
		14'h1092: color = 2'b11;
		14'h1093: color = 2'b11;
		14'h1094: color = 2'b11;
		14'h1095: color = 2'b11;
		14'h1096: color = 2'b11;
		14'h1097: color = 2'b11;
		14'h1098: color = 2'b11;
		14'h1099: color = 2'b11;
		14'h109a: color = 2'b11;
		14'h109b: color = 2'b11;
		14'h109c: color = 2'b11;
		14'h109d: color = 2'b11;
		14'h109e: color = 2'b11;
		14'h109f: color = 2'b11;
		14'h10a0: color = 2'b11;
		14'h10a1: color = 2'b11;
		14'h10a2: color = 2'b11;
		14'h10a3: color = 2'b01;
		14'h10a4: color = 2'b00;
		14'h10a5: color = 2'b00;
		14'h10a6: color = 2'b00;
		14'h10a7: color = 2'b00;
		14'h10a8: color = 2'b00;
		14'h10a9: color = 2'b00;
		14'h10aa: color = 2'b01;
		14'h10ab: color = 2'b01;
		14'h10ac: color = 2'b00;
		14'h10ad: color = 2'b01;
		14'h10ae: color = 2'b00;
		14'h10af: color = 2'b01;
		14'h10b0: color = 2'b00;
		14'h10b1: color = 2'b00;
		14'h10b2: color = 2'b00;
		14'h10b3: color = 2'b00;
		14'h10b4: color = 2'b00;
		14'h10b5: color = 2'b00;
		14'h10b6: color = 2'b00;
		14'h10b7: color = 2'b01;
		14'h10b8: color = 2'b01;
		14'h10b9: color = 2'b01;
		14'h10ba: color = 2'b01;
		14'h10bb: color = 2'b00;
		14'h10bc: color = 2'b01;
		14'h10bd: color = 2'b00;
		14'h10be: color = 2'b00;
		14'h10bf: color = 2'b00;
		14'h10c0: color = 2'b01;
		14'h10c1: color = 2'b00;
		14'h10c2: color = 2'b00;
		14'h10c3: color = 2'b00;
		14'h10c4: color = 2'b00;
		14'h10c5: color = 2'b00;
		14'h10c6: color = 2'b00;
		14'h10c7: color = 2'b00;
		14'h10c8: color = 2'b00;
		14'h10c9: color = 2'b00;
		14'h10ca: color = 2'b00;
		14'h10cb: color = 2'b00;
		14'h10cc: color = 2'b00;
		14'h10cd: color = 2'b00;
		14'h10ce: color = 2'b00;
		14'h10cf: color = 2'b00;
		14'h10d0: color = 2'b00;
		14'h10d1: color = 2'b00;
		14'h10d2: color = 2'b00;
		14'h10d3: color = 2'b01;
		14'h10d4: color = 2'b01;
		14'h10d5: color = 2'b01;
		14'h10d6: color = 2'b01;
		14'h10d7: color = 2'b01;
		14'h10d8: color = 2'b01;
		14'h10d9: color = 2'b01;
		14'h10da: color = 2'b01;
		14'h10db: color = 2'b01;
		14'h10dc: color = 2'b10;
		14'h10dd: color = 2'b01;
		14'h10de: color = 2'b01;
		14'h10df: color = 2'b00;
		14'h10e0: color = 2'b00;
		14'h10e1: color = 2'b00;
		14'h10e2: color = 2'b00;
		14'h10e3: color = 2'b00;
		14'h10e4: color = 2'b00;
		14'h10e5: color = 2'b00;
		14'h10e6: color = 2'b00;
		14'h10e7: color = 2'b01;
		14'h10e8: color = 2'b01;
		14'h10e9: color = 2'b11;
		14'h10ea: color = 2'b11;
		14'h10eb: color = 2'b11;
		14'h10ec: color = 2'b11;
		14'h10ed: color = 2'b11;
		14'h10ee: color = 2'b11;
		14'h10ef: color = 2'b11;
		14'h10f0: color = 2'b11;
		14'h10f1: color = 2'b11;
		14'h10f2: color = 2'b11;
		14'h10f3: color = 2'b11;
		14'h10f4: color = 2'b11;
		14'h10f5: color = 2'b11;
		14'h10f6: color = 2'b11;
		14'h10f7: color = 2'b11;
		14'h10f8: color = 2'b11;
		14'h10f9: color = 2'b11;
		14'h10fa: color = 2'b11;
		14'h10fb: color = 2'b11;
		14'h10fc: color = 2'b11;
		14'h10fd: color = 2'b11;
		14'h10fe: color = 2'b11;
		14'h10ff: color = 2'b11;
		14'h1100: color = 2'b11;
		14'h1101: color = 2'b11;
		14'h1102: color = 2'b11;
		14'h1103: color = 2'b11;
		14'h1104: color = 2'b11;
		14'h1105: color = 2'b11;
		14'h1106: color = 2'b11;
		14'h1107: color = 2'b11;
		14'h1108: color = 2'b11;
		14'h1109: color = 2'b11;
		14'h110a: color = 2'b11;
		14'h110b: color = 2'b11;
		14'h110c: color = 2'b11;
		14'h110d: color = 2'b11;
		14'h110e: color = 2'b11;
		14'h110f: color = 2'b11;
		14'h1110: color = 2'b11;
		14'h1111: color = 2'b11;
		14'h1112: color = 2'b11;
		14'h1113: color = 2'b11;
		14'h1114: color = 2'b11;
		14'h1115: color = 2'b11;
		14'h1116: color = 2'b11;
		14'h1117: color = 2'b11;
		14'h1118: color = 2'b11;
		14'h1119: color = 2'b11;
		14'h111a: color = 2'b11;
		14'h111b: color = 2'b11;
		14'h111c: color = 2'b11;
		14'h111d: color = 2'b11;
		14'h111e: color = 2'b11;
		14'h111f: color = 2'b11;
		14'h1120: color = 2'b11;
		14'h1121: color = 2'b11;
		14'h1122: color = 2'b10;
		14'h1123: color = 2'b00;
		14'h1124: color = 2'b00;
		14'h1125: color = 2'b00;
		14'h1126: color = 2'b00;
		14'h1127: color = 2'b00;
		14'h1128: color = 2'b00;
		14'h1129: color = 2'b01;
		14'h112a: color = 2'b00;
		14'h112b: color = 2'b00;
		14'h112c: color = 2'b01;
		14'h112d: color = 2'b00;
		14'h112e: color = 2'b01;
		14'h112f: color = 2'b00;
		14'h1130: color = 2'b00;
		14'h1131: color = 2'b00;
		14'h1132: color = 2'b00;
		14'h1133: color = 2'b00;
		14'h1134: color = 2'b00;
		14'h1135: color = 2'b00;
		14'h1136: color = 2'b00;
		14'h1137: color = 2'b00;
		14'h1138: color = 2'b00;
		14'h1139: color = 2'b00;
		14'h113a: color = 2'b01;
		14'h113b: color = 2'b01;
		14'h113c: color = 2'b01;
		14'h113d: color = 2'b00;
		14'h113e: color = 2'b00;
		14'h113f: color = 2'b00;
		14'h1140: color = 2'b00;
		14'h1141: color = 2'b00;
		14'h1142: color = 2'b00;
		14'h1143: color = 2'b00;
		14'h1144: color = 2'b00;
		14'h1145: color = 2'b00;
		14'h1146: color = 2'b00;
		14'h1147: color = 2'b00;
		14'h1148: color = 2'b00;
		14'h1149: color = 2'b00;
		14'h114a: color = 2'b00;
		14'h114b: color = 2'b00;
		14'h114c: color = 2'b00;
		14'h114d: color = 2'b00;
		14'h114e: color = 2'b00;
		14'h114f: color = 2'b01;
		14'h1150: color = 2'b00;
		14'h1151: color = 2'b00;
		14'h1152: color = 2'b00;
		14'h1153: color = 2'b01;
		14'h1154: color = 2'b00;
		14'h1155: color = 2'b01;
		14'h1156: color = 2'b01;
		14'h1157: color = 2'b01;
		14'h1158: color = 2'b01;
		14'h1159: color = 2'b01;
		14'h115a: color = 2'b01;
		14'h115b: color = 2'b10;
		14'h115c: color = 2'b01;
		14'h115d: color = 2'b10;
		14'h115e: color = 2'b01;
		14'h115f: color = 2'b00;
		14'h1160: color = 2'b00;
		14'h1161: color = 2'b00;
		14'h1162: color = 2'b00;
		14'h1163: color = 2'b00;
		14'h1164: color = 2'b00;
		14'h1165: color = 2'b00;
		14'h1166: color = 2'b00;
		14'h1167: color = 2'b01;
		14'h1168: color = 2'b01;
		14'h1169: color = 2'b11;
		14'h116a: color = 2'b11;
		14'h116b: color = 2'b11;
		14'h116c: color = 2'b11;
		14'h116d: color = 2'b11;
		14'h116e: color = 2'b11;
		14'h116f: color = 2'b11;
		14'h1170: color = 2'b11;
		14'h1171: color = 2'b11;
		14'h1172: color = 2'b11;
		14'h1173: color = 2'b11;
		14'h1174: color = 2'b11;
		14'h1175: color = 2'b11;
		14'h1176: color = 2'b11;
		14'h1177: color = 2'b11;
		14'h1178: color = 2'b11;
		14'h1179: color = 2'b11;
		14'h117a: color = 2'b11;
		14'h117b: color = 2'b11;
		14'h117c: color = 2'b11;
		14'h117d: color = 2'b11;
		14'h117e: color = 2'b11;
		14'h117f: color = 2'b11;
		14'h1180: color = 2'b11;
		14'h1181: color = 2'b11;
		14'h1182: color = 2'b11;
		14'h1183: color = 2'b11;
		14'h1184: color = 2'b11;
		14'h1185: color = 2'b11;
		14'h1186: color = 2'b11;
		14'h1187: color = 2'b11;
		14'h1188: color = 2'b11;
		14'h1189: color = 2'b11;
		14'h118a: color = 2'b11;
		14'h118b: color = 2'b11;
		14'h118c: color = 2'b11;
		14'h118d: color = 2'b11;
		14'h118e: color = 2'b11;
		14'h118f: color = 2'b11;
		14'h1190: color = 2'b11;
		14'h1191: color = 2'b11;
		14'h1192: color = 2'b11;
		14'h1193: color = 2'b11;
		14'h1194: color = 2'b11;
		14'h1195: color = 2'b11;
		14'h1196: color = 2'b11;
		14'h1197: color = 2'b11;
		14'h1198: color = 2'b11;
		14'h1199: color = 2'b11;
		14'h119a: color = 2'b11;
		14'h119b: color = 2'b11;
		14'h119c: color = 2'b11;
		14'h119d: color = 2'b11;
		14'h119e: color = 2'b11;
		14'h119f: color = 2'b11;
		14'h11a0: color = 2'b11;
		14'h11a1: color = 2'b10;
		14'h11a2: color = 2'b01;
		14'h11a3: color = 2'b01;
		14'h11a4: color = 2'b00;
		14'h11a5: color = 2'b00;
		14'h11a6: color = 2'b00;
		14'h11a7: color = 2'b01;
		14'h11a8: color = 2'b01;
		14'h11a9: color = 2'b00;
		14'h11aa: color = 2'b01;
		14'h11ab: color = 2'b01;
		14'h11ac: color = 2'b00;
		14'h11ad: color = 2'b01;
		14'h11ae: color = 2'b01;
		14'h11af: color = 2'b00;
		14'h11b0: color = 2'b01;
		14'h11b1: color = 2'b00;
		14'h11b2: color = 2'b00;
		14'h11b3: color = 2'b00;
		14'h11b4: color = 2'b00;
		14'h11b5: color = 2'b00;
		14'h11b6: color = 2'b00;
		14'h11b7: color = 2'b01;
		14'h11b8: color = 2'b01;
		14'h11b9: color = 2'b01;
		14'h11ba: color = 2'b01;
		14'h11bb: color = 2'b01;
		14'h11bc: color = 2'b00;
		14'h11bd: color = 2'b00;
		14'h11be: color = 2'b00;
		14'h11bf: color = 2'b01;
		14'h11c0: color = 2'b00;
		14'h11c1: color = 2'b00;
		14'h11c2: color = 2'b00;
		14'h11c3: color = 2'b00;
		14'h11c4: color = 2'b01;
		14'h11c5: color = 2'b00;
		14'h11c6: color = 2'b00;
		14'h11c7: color = 2'b00;
		14'h11c8: color = 2'b00;
		14'h11c9: color = 2'b00;
		14'h11ca: color = 2'b00;
		14'h11cb: color = 2'b01;
		14'h11cc: color = 2'b00;
		14'h11cd: color = 2'b01;
		14'h11ce: color = 2'b01;
		14'h11cf: color = 2'b01;
		14'h11d0: color = 2'b01;
		14'h11d1: color = 2'b01;
		14'h11d2: color = 2'b01;
		14'h11d3: color = 2'b01;
		14'h11d4: color = 2'b01;
		14'h11d5: color = 2'b01;
		14'h11d6: color = 2'b10;
		14'h11d7: color = 2'b01;
		14'h11d8: color = 2'b01;
		14'h11d9: color = 2'b10;
		14'h11da: color = 2'b10;
		14'h11db: color = 2'b01;
		14'h11dc: color = 2'b10;
		14'h11dd: color = 2'b10;
		14'h11de: color = 2'b01;
		14'h11df: color = 2'b01;
		14'h11e0: color = 2'b00;
		14'h11e1: color = 2'b00;
		14'h11e2: color = 2'b00;
		14'h11e3: color = 2'b00;
		14'h11e4: color = 2'b00;
		14'h11e5: color = 2'b00;
		14'h11e6: color = 2'b00;
		14'h11e7: color = 2'b00;
		14'h11e8: color = 2'b00;
		14'h11e9: color = 2'b11;
		14'h11ea: color = 2'b11;
		14'h11eb: color = 2'b11;
		14'h11ec: color = 2'b11;
		14'h11ed: color = 2'b11;
		14'h11ee: color = 2'b11;
		14'h11ef: color = 2'b11;
		14'h11f0: color = 2'b11;
		14'h11f1: color = 2'b11;
		14'h11f2: color = 2'b11;
		14'h11f3: color = 2'b11;
		14'h11f4: color = 2'b11;
		14'h11f5: color = 2'b11;
		14'h11f6: color = 2'b11;
		14'h11f7: color = 2'b11;
		14'h11f8: color = 2'b11;
		14'h11f9: color = 2'b11;
		14'h11fa: color = 2'b11;
		14'h11fb: color = 2'b11;
		14'h11fc: color = 2'b11;
		14'h11fd: color = 2'b11;
		14'h11fe: color = 2'b11;
		14'h11ff: color = 2'b11;
		14'h1200: color = 2'b11;
		14'h1201: color = 2'b11;
		14'h1202: color = 2'b11;
		14'h1203: color = 2'b11;
		14'h1204: color = 2'b11;
		14'h1205: color = 2'b11;
		14'h1206: color = 2'b11;
		14'h1207: color = 2'b11;
		14'h1208: color = 2'b11;
		14'h1209: color = 2'b11;
		14'h120a: color = 2'b11;
		14'h120b: color = 2'b11;
		14'h120c: color = 2'b11;
		14'h120d: color = 2'b11;
		14'h120e: color = 2'b11;
		14'h120f: color = 2'b11;
		14'h1210: color = 2'b11;
		14'h1211: color = 2'b11;
		14'h1212: color = 2'b11;
		14'h1213: color = 2'b11;
		14'h1214: color = 2'b11;
		14'h1215: color = 2'b11;
		14'h1216: color = 2'b11;
		14'h1217: color = 2'b11;
		14'h1218: color = 2'b11;
		14'h1219: color = 2'b11;
		14'h121a: color = 2'b11;
		14'h121b: color = 2'b11;
		14'h121c: color = 2'b11;
		14'h121d: color = 2'b11;
		14'h121e: color = 2'b11;
		14'h121f: color = 2'b11;
		14'h1220: color = 2'b11;
		14'h1221: color = 2'b10;
		14'h1222: color = 2'b01;
		14'h1223: color = 2'b00;
		14'h1224: color = 2'b01;
		14'h1225: color = 2'b00;
		14'h1226: color = 2'b00;
		14'h1227: color = 2'b00;
		14'h1228: color = 2'b00;
		14'h1229: color = 2'b00;
		14'h122a: color = 2'b01;
		14'h122b: color = 2'b00;
		14'h122c: color = 2'b01;
		14'h122d: color = 2'b00;
		14'h122e: color = 2'b01;
		14'h122f: color = 2'b00;
		14'h1230: color = 2'b00;
		14'h1231: color = 2'b00;
		14'h1232: color = 2'b00;
		14'h1233: color = 2'b00;
		14'h1234: color = 2'b00;
		14'h1235: color = 2'b00;
		14'h1236: color = 2'b00;
		14'h1237: color = 2'b01;
		14'h1238: color = 2'b01;
		14'h1239: color = 2'b00;
		14'h123a: color = 2'b01;
		14'h123b: color = 2'b00;
		14'h123c: color = 2'b00;
		14'h123d: color = 2'b01;
		14'h123e: color = 2'b00;
		14'h123f: color = 2'b00;
		14'h1240: color = 2'b00;
		14'h1241: color = 2'b00;
		14'h1242: color = 2'b00;
		14'h1243: color = 2'b00;
		14'h1244: color = 2'b00;
		14'h1245: color = 2'b01;
		14'h1246: color = 2'b00;
		14'h1247: color = 2'b00;
		14'h1248: color = 2'b00;
		14'h1249: color = 2'b01;
		14'h124a: color = 2'b00;
		14'h124b: color = 2'b01;
		14'h124c: color = 2'b01;
		14'h124d: color = 2'b00;
		14'h124e: color = 2'b01;
		14'h124f: color = 2'b01;
		14'h1250: color = 2'b01;
		14'h1251: color = 2'b01;
		14'h1252: color = 2'b10;
		14'h1253: color = 2'b01;
		14'h1254: color = 2'b10;
		14'h1255: color = 2'b10;
		14'h1256: color = 2'b01;
		14'h1257: color = 2'b10;
		14'h1258: color = 2'b10;
		14'h1259: color = 2'b01;
		14'h125a: color = 2'b10;
		14'h125b: color = 2'b10;
		14'h125c: color = 2'b10;
		14'h125d: color = 2'b01;
		14'h125e: color = 2'b10;
		14'h125f: color = 2'b01;
		14'h1260: color = 2'b00;
		14'h1261: color = 2'b00;
		14'h1262: color = 2'b00;
		14'h1263: color = 2'b00;
		14'h1264: color = 2'b00;
		14'h1265: color = 2'b00;
		14'h1266: color = 2'b00;
		14'h1267: color = 2'b00;
		14'h1268: color = 2'b00;
		14'h1269: color = 2'b00;
		14'h126a: color = 2'b10;
		14'h126b: color = 2'b11;
		14'h126c: color = 2'b11;
		14'h126d: color = 2'b11;
		14'h126e: color = 2'b11;
		14'h126f: color = 2'b11;
		14'h1270: color = 2'b11;
		14'h1271: color = 2'b11;
		14'h1272: color = 2'b11;
		14'h1273: color = 2'b11;
		14'h1274: color = 2'b11;
		14'h1275: color = 2'b11;
		14'h1276: color = 2'b11;
		14'h1277: color = 2'b11;
		14'h1278: color = 2'b11;
		14'h1279: color = 2'b11;
		14'h127a: color = 2'b11;
		14'h127b: color = 2'b11;
		14'h127c: color = 2'b11;
		14'h127d: color = 2'b11;
		14'h127e: color = 2'b11;
		14'h127f: color = 2'b11;
		14'h1280: color = 2'b11;
		14'h1281: color = 2'b11;
		14'h1282: color = 2'b11;
		14'h1283: color = 2'b11;
		14'h1284: color = 2'b11;
		14'h1285: color = 2'b11;
		14'h1286: color = 2'b11;
		14'h1287: color = 2'b11;
		14'h1288: color = 2'b11;
		14'h1289: color = 2'b11;
		14'h128a: color = 2'b11;
		14'h128b: color = 2'b11;
		14'h128c: color = 2'b11;
		14'h128d: color = 2'b11;
		14'h128e: color = 2'b11;
		14'h128f: color = 2'b11;
		14'h1290: color = 2'b11;
		14'h1291: color = 2'b11;
		14'h1292: color = 2'b11;
		14'h1293: color = 2'b11;
		14'h1294: color = 2'b11;
		14'h1295: color = 2'b11;
		14'h1296: color = 2'b11;
		14'h1297: color = 2'b11;
		14'h1298: color = 2'b11;
		14'h1299: color = 2'b11;
		14'h129a: color = 2'b11;
		14'h129b: color = 2'b11;
		14'h129c: color = 2'b11;
		14'h129d: color = 2'b11;
		14'h129e: color = 2'b11;
		14'h129f: color = 2'b11;
		14'h12a0: color = 2'b11;
		14'h12a1: color = 2'b10;
		14'h12a2: color = 2'b00;
		14'h12a3: color = 2'b01;
		14'h12a4: color = 2'b01;
		14'h12a5: color = 2'b00;
		14'h12a6: color = 2'b00;
		14'h12a7: color = 2'b01;
		14'h12a8: color = 2'b01;
		14'h12a9: color = 2'b00;
		14'h12aa: color = 2'b01;
		14'h12ab: color = 2'b00;
		14'h12ac: color = 2'b00;
		14'h12ad: color = 2'b00;
		14'h12ae: color = 2'b01;
		14'h12af: color = 2'b00;
		14'h12b0: color = 2'b00;
		14'h12b1: color = 2'b00;
		14'h12b2: color = 2'b00;
		14'h12b3: color = 2'b00;
		14'h12b4: color = 2'b00;
		14'h12b5: color = 2'b01;
		14'h12b6: color = 2'b01;
		14'h12b7: color = 2'b01;
		14'h12b8: color = 2'b01;
		14'h12b9: color = 2'b01;
		14'h12ba: color = 2'b01;
		14'h12bb: color = 2'b00;
		14'h12bc: color = 2'b01;
		14'h12bd: color = 2'b00;
		14'h12be: color = 2'b00;
		14'h12bf: color = 2'b01;
		14'h12c0: color = 2'b00;
		14'h12c1: color = 2'b00;
		14'h12c2: color = 2'b00;
		14'h12c3: color = 2'b00;
		14'h12c4: color = 2'b01;
		14'h12c5: color = 2'b01;
		14'h12c6: color = 2'b01;
		14'h12c7: color = 2'b01;
		14'h12c8: color = 2'b01;
		14'h12c9: color = 2'b01;
		14'h12ca: color = 2'b01;
		14'h12cb: color = 2'b01;
		14'h12cc: color = 2'b01;
		14'h12cd: color = 2'b10;
		14'h12ce: color = 2'b01;
		14'h12cf: color = 2'b01;
		14'h12d0: color = 2'b01;
		14'h12d1: color = 2'b10;
		14'h12d2: color = 2'b01;
		14'h12d3: color = 2'b10;
		14'h12d4: color = 2'b10;
		14'h12d5: color = 2'b10;
		14'h12d6: color = 2'b10;
		14'h12d7: color = 2'b10;
		14'h12d8: color = 2'b10;
		14'h12d9: color = 2'b10;
		14'h12da: color = 2'b10;
		14'h12db: color = 2'b01;
		14'h12dc: color = 2'b10;
		14'h12dd: color = 2'b01;
		14'h12de: color = 2'b10;
		14'h12df: color = 2'b01;
		14'h12e0: color = 2'b00;
		14'h12e1: color = 2'b00;
		14'h12e2: color = 2'b00;
		14'h12e3: color = 2'b00;
		14'h12e4: color = 2'b00;
		14'h12e5: color = 2'b00;
		14'h12e6: color = 2'b00;
		14'h12e7: color = 2'b00;
		14'h12e8: color = 2'b00;
		14'h12e9: color = 2'b00;
		14'h12ea: color = 2'b00;
		14'h12eb: color = 2'b11;
		14'h12ec: color = 2'b11;
		14'h12ed: color = 2'b11;
		14'h12ee: color = 2'b11;
		14'h12ef: color = 2'b11;
		14'h12f0: color = 2'b11;
		14'h12f1: color = 2'b11;
		14'h12f2: color = 2'b11;
		14'h12f3: color = 2'b11;
		14'h12f4: color = 2'b11;
		14'h12f5: color = 2'b11;
		14'h12f6: color = 2'b11;
		14'h12f7: color = 2'b11;
		14'h12f8: color = 2'b11;
		14'h12f9: color = 2'b11;
		14'h12fa: color = 2'b11;
		14'h12fb: color = 2'b11;
		14'h12fc: color = 2'b11;
		14'h12fd: color = 2'b11;
		14'h12fe: color = 2'b11;
		14'h12ff: color = 2'b11;
		14'h1300: color = 2'b11;
		14'h1301: color = 2'b11;
		14'h1302: color = 2'b11;
		14'h1303: color = 2'b11;
		14'h1304: color = 2'b11;
		14'h1305: color = 2'b11;
		14'h1306: color = 2'b11;
		14'h1307: color = 2'b11;
		14'h1308: color = 2'b11;
		14'h1309: color = 2'b11;
		14'h130a: color = 2'b11;
		14'h130b: color = 2'b11;
		14'h130c: color = 2'b11;
		14'h130d: color = 2'b11;
		14'h130e: color = 2'b11;
		14'h130f: color = 2'b11;
		14'h1310: color = 2'b11;
		14'h1311: color = 2'b11;
		14'h1312: color = 2'b11;
		14'h1313: color = 2'b11;
		14'h1314: color = 2'b11;
		14'h1315: color = 2'b11;
		14'h1316: color = 2'b11;
		14'h1317: color = 2'b11;
		14'h1318: color = 2'b11;
		14'h1319: color = 2'b11;
		14'h131a: color = 2'b11;
		14'h131b: color = 2'b11;
		14'h131c: color = 2'b11;
		14'h131d: color = 2'b11;
		14'h131e: color = 2'b11;
		14'h131f: color = 2'b11;
		14'h1320: color = 2'b11;
		14'h1321: color = 2'b10;
		14'h1322: color = 2'b00;
		14'h1323: color = 2'b01;
		14'h1324: color = 2'b00;
		14'h1325: color = 2'b01;
		14'h1326: color = 2'b00;
		14'h1327: color = 2'b00;
		14'h1328: color = 2'b00;
		14'h1329: color = 2'b00;
		14'h132a: color = 2'b00;
		14'h132b: color = 2'b01;
		14'h132c: color = 2'b00;
		14'h132d: color = 2'b00;
		14'h132e: color = 2'b00;
		14'h132f: color = 2'b00;
		14'h1330: color = 2'b01;
		14'h1331: color = 2'b01;
		14'h1332: color = 2'b00;
		14'h1333: color = 2'b00;
		14'h1334: color = 2'b00;
		14'h1335: color = 2'b00;
		14'h1336: color = 2'b10;
		14'h1337: color = 2'b10;
		14'h1338: color = 2'b10;
		14'h1339: color = 2'b11;
		14'h133a: color = 2'b11;
		14'h133b: color = 2'b11;
		14'h133c: color = 2'b10;
		14'h133d: color = 2'b10;
		14'h133e: color = 2'b01;
		14'h133f: color = 2'b01;
		14'h1340: color = 2'b00;
		14'h1341: color = 2'b01;
		14'h1342: color = 2'b01;
		14'h1343: color = 2'b01;
		14'h1344: color = 2'b01;
		14'h1345: color = 2'b01;
		14'h1346: color = 2'b10;
		14'h1347: color = 2'b10;
		14'h1348: color = 2'b10;
		14'h1349: color = 2'b10;
		14'h134a: color = 2'b10;
		14'h134b: color = 2'b10;
		14'h134c: color = 2'b10;
		14'h134d: color = 2'b10;
		14'h134e: color = 2'b10;
		14'h134f: color = 2'b10;
		14'h1350: color = 2'b10;
		14'h1351: color = 2'b10;
		14'h1352: color = 2'b10;
		14'h1353: color = 2'b10;
		14'h1354: color = 2'b10;
		14'h1355: color = 2'b10;
		14'h1356: color = 2'b10;
		14'h1357: color = 2'b01;
		14'h1358: color = 2'b01;
		14'h1359: color = 2'b10;
		14'h135a: color = 2'b10;
		14'h135b: color = 2'b10;
		14'h135c: color = 2'b10;
		14'h135d: color = 2'b10;
		14'h135e: color = 2'b10;
		14'h135f: color = 2'b01;
		14'h1360: color = 2'b00;
		14'h1361: color = 2'b00;
		14'h1362: color = 2'b00;
		14'h1363: color = 2'b00;
		14'h1364: color = 2'b00;
		14'h1365: color = 2'b00;
		14'h1366: color = 2'b00;
		14'h1367: color = 2'b00;
		14'h1368: color = 2'b00;
		14'h1369: color = 2'b00;
		14'h136a: color = 2'b00;
		14'h136b: color = 2'b11;
		14'h136c: color = 2'b11;
		14'h136d: color = 2'b11;
		14'h136e: color = 2'b11;
		14'h136f: color = 2'b11;
		14'h1370: color = 2'b11;
		14'h1371: color = 2'b11;
		14'h1372: color = 2'b11;
		14'h1373: color = 2'b11;
		14'h1374: color = 2'b11;
		14'h1375: color = 2'b11;
		14'h1376: color = 2'b11;
		14'h1377: color = 2'b11;
		14'h1378: color = 2'b11;
		14'h1379: color = 2'b11;
		14'h137a: color = 2'b11;
		14'h137b: color = 2'b11;
		14'h137c: color = 2'b11;
		14'h137d: color = 2'b11;
		14'h137e: color = 2'b11;
		14'h137f: color = 2'b11;
		14'h1380: color = 2'b11;
		14'h1381: color = 2'b11;
		14'h1382: color = 2'b11;
		14'h1383: color = 2'b11;
		14'h1384: color = 2'b11;
		14'h1385: color = 2'b11;
		14'h1386: color = 2'b11;
		14'h1387: color = 2'b11;
		14'h1388: color = 2'b11;
		14'h1389: color = 2'b11;
		14'h138a: color = 2'b11;
		14'h138b: color = 2'b11;
		14'h138c: color = 2'b11;
		14'h138d: color = 2'b11;
		14'h138e: color = 2'b11;
		14'h138f: color = 2'b11;
		14'h1390: color = 2'b11;
		14'h1391: color = 2'b11;
		14'h1392: color = 2'b11;
		14'h1393: color = 2'b11;
		14'h1394: color = 2'b11;
		14'h1395: color = 2'b11;
		14'h1396: color = 2'b11;
		14'h1397: color = 2'b11;
		14'h1398: color = 2'b11;
		14'h1399: color = 2'b11;
		14'h139a: color = 2'b11;
		14'h139b: color = 2'b11;
		14'h139c: color = 2'b11;
		14'h139d: color = 2'b11;
		14'h139e: color = 2'b11;
		14'h139f: color = 2'b11;
		14'h13a0: color = 2'b11;
		14'h13a1: color = 2'b10;
		14'h13a2: color = 2'b00;
		14'h13a3: color = 2'b00;
		14'h13a4: color = 2'b00;
		14'h13a5: color = 2'b01;
		14'h13a6: color = 2'b00;
		14'h13a7: color = 2'b01;
		14'h13a8: color = 2'b01;
		14'h13a9: color = 2'b00;
		14'h13aa: color = 2'b01;
		14'h13ab: color = 2'b00;
		14'h13ac: color = 2'b01;
		14'h13ad: color = 2'b00;
		14'h13ae: color = 2'b00;
		14'h13af: color = 2'b00;
		14'h13b0: color = 2'b01;
		14'h13b1: color = 2'b00;
		14'h13b2: color = 2'b01;
		14'h13b3: color = 2'b00;
		14'h13b4: color = 2'b00;
		14'h13b5: color = 2'b01;
		14'h13b6: color = 2'b10;
		14'h13b7: color = 2'b11;
		14'h13b8: color = 2'b11;
		14'h13b9: color = 2'b11;
		14'h13ba: color = 2'b11;
		14'h13bb: color = 2'b11;
		14'h13bc: color = 2'b11;
		14'h13bd: color = 2'b11;
		14'h13be: color = 2'b11;
		14'h13bf: color = 2'b10;
		14'h13c0: color = 2'b11;
		14'h13c1: color = 2'b10;
		14'h13c2: color = 2'b10;
		14'h13c3: color = 2'b11;
		14'h13c4: color = 2'b10;
		14'h13c5: color = 2'b10;
		14'h13c6: color = 2'b10;
		14'h13c7: color = 2'b10;
		14'h13c8: color = 2'b10;
		14'h13c9: color = 2'b10;
		14'h13ca: color = 2'b10;
		14'h13cb: color = 2'b10;
		14'h13cc: color = 2'b10;
		14'h13cd: color = 2'b10;
		14'h13ce: color = 2'b10;
		14'h13cf: color = 2'b10;
		14'h13d0: color = 2'b10;
		14'h13d1: color = 2'b10;
		14'h13d2: color = 2'b10;
		14'h13d3: color = 2'b10;
		14'h13d4: color = 2'b10;
		14'h13d5: color = 2'b10;
		14'h13d6: color = 2'b10;
		14'h13d7: color = 2'b10;
		14'h13d8: color = 2'b10;
		14'h13d9: color = 2'b10;
		14'h13da: color = 2'b10;
		14'h13db: color = 2'b01;
		14'h13dc: color = 2'b10;
		14'h13dd: color = 2'b01;
		14'h13de: color = 2'b10;
		14'h13df: color = 2'b01;
		14'h13e0: color = 2'b00;
		14'h13e1: color = 2'b00;
		14'h13e2: color = 2'b00;
		14'h13e3: color = 2'b00;
		14'h13e4: color = 2'b00;
		14'h13e5: color = 2'b00;
		14'h13e6: color = 2'b00;
		14'h13e7: color = 2'b00;
		14'h13e8: color = 2'b00;
		14'h13e9: color = 2'b00;
		14'h13ea: color = 2'b00;
		14'h13eb: color = 2'b11;
		14'h13ec: color = 2'b11;
		14'h13ed: color = 2'b11;
		14'h13ee: color = 2'b11;
		14'h13ef: color = 2'b11;
		14'h13f0: color = 2'b11;
		14'h13f1: color = 2'b11;
		14'h13f2: color = 2'b11;
		14'h13f3: color = 2'b11;
		14'h13f4: color = 2'b11;
		14'h13f5: color = 2'b11;
		14'h13f6: color = 2'b11;
		14'h13f7: color = 2'b11;
		14'h13f8: color = 2'b11;
		14'h13f9: color = 2'b11;
		14'h13fa: color = 2'b11;
		14'h13fb: color = 2'b11;
		14'h13fc: color = 2'b11;
		14'h13fd: color = 2'b11;
		14'h13fe: color = 2'b11;
		14'h13ff: color = 2'b11;
		14'h1400: color = 2'b11;
		14'h1401: color = 2'b11;
		14'h1402: color = 2'b11;
		14'h1403: color = 2'b11;
		14'h1404: color = 2'b11;
		14'h1405: color = 2'b11;
		14'h1406: color = 2'b11;
		14'h1407: color = 2'b11;
		14'h1408: color = 2'b11;
		14'h1409: color = 2'b11;
		14'h140a: color = 2'b11;
		14'h140b: color = 2'b11;
		14'h140c: color = 2'b11;
		14'h140d: color = 2'b11;
		14'h140e: color = 2'b11;
		14'h140f: color = 2'b11;
		14'h1410: color = 2'b11;
		14'h1411: color = 2'b11;
		14'h1412: color = 2'b11;
		14'h1413: color = 2'b11;
		14'h1414: color = 2'b11;
		14'h1415: color = 2'b11;
		14'h1416: color = 2'b11;
		14'h1417: color = 2'b11;
		14'h1418: color = 2'b11;
		14'h1419: color = 2'b11;
		14'h141a: color = 2'b11;
		14'h141b: color = 2'b11;
		14'h141c: color = 2'b11;
		14'h141d: color = 2'b11;
		14'h141e: color = 2'b11;
		14'h141f: color = 2'b11;
		14'h1420: color = 2'b11;
		14'h1421: color = 2'b10;
		14'h1422: color = 2'b00;
		14'h1423: color = 2'b00;
		14'h1424: color = 2'b00;
		14'h1425: color = 2'b01;
		14'h1426: color = 2'b00;
		14'h1427: color = 2'b01;
		14'h1428: color = 2'b01;
		14'h1429: color = 2'b00;
		14'h142a: color = 2'b01;
		14'h142b: color = 2'b00;
		14'h142c: color = 2'b01;
		14'h142d: color = 2'b00;
		14'h142e: color = 2'b00;
		14'h142f: color = 2'b00;
		14'h1430: color = 2'b01;
		14'h1431: color = 2'b00;
		14'h1432: color = 2'b01;
		14'h1433: color = 2'b00;
		14'h1434: color = 2'b00;
		14'h1435: color = 2'b01;
		14'h1436: color = 2'b10;
		14'h1437: color = 2'b11;
		14'h1438: color = 2'b11;
		14'h1439: color = 2'b11;
		14'h143a: color = 2'b11;
		14'h143b: color = 2'b11;
		14'h143c: color = 2'b11;
		14'h143d: color = 2'b11;
		14'h143e: color = 2'b11;
		14'h143f: color = 2'b10;
		14'h1440: color = 2'b11;
		14'h1441: color = 2'b10;
		14'h1442: color = 2'b10;
		14'h1443: color = 2'b11;
		14'h1444: color = 2'b10;
		14'h1445: color = 2'b10;
		14'h1446: color = 2'b10;
		14'h1447: color = 2'b10;
		14'h1448: color = 2'b10;
		14'h1449: color = 2'b10;
		14'h144a: color = 2'b10;
		14'h144b: color = 2'b10;
		14'h144c: color = 2'b10;
		14'h144d: color = 2'b10;
		14'h144e: color = 2'b10;
		14'h144f: color = 2'b10;
		14'h1450: color = 2'b10;
		14'h1451: color = 2'b10;
		14'h1452: color = 2'b10;
		14'h1453: color = 2'b10;
		14'h1454: color = 2'b10;
		14'h1455: color = 2'b10;
		14'h1456: color = 2'b10;
		14'h1457: color = 2'b10;
		14'h1458: color = 2'b10;
		14'h1459: color = 2'b10;
		14'h145a: color = 2'b10;
		14'h145b: color = 2'b01;
		14'h145c: color = 2'b10;
		14'h145d: color = 2'b01;
		14'h145e: color = 2'b10;
		14'h145f: color = 2'b01;
		14'h1460: color = 2'b00;
		14'h1461: color = 2'b00;
		14'h1462: color = 2'b00;
		14'h1463: color = 2'b00;
		14'h1464: color = 2'b00;
		14'h1465: color = 2'b00;
		14'h1466: color = 2'b00;
		14'h1467: color = 2'b00;
		14'h1468: color = 2'b00;
		14'h1469: color = 2'b00;
		14'h146a: color = 2'b00;
		14'h146b: color = 2'b11;
		14'h146c: color = 2'b11;
		14'h146d: color = 2'b11;
		14'h146e: color = 2'b11;
		14'h146f: color = 2'b11;
		14'h1470: color = 2'b11;
		14'h1471: color = 2'b11;
		14'h1472: color = 2'b11;
		14'h1473: color = 2'b11;
		14'h1474: color = 2'b11;
		14'h1475: color = 2'b11;
		14'h1476: color = 2'b11;
		14'h1477: color = 2'b11;
		14'h1478: color = 2'b11;
		14'h1479: color = 2'b11;
		14'h147a: color = 2'b11;
		14'h147b: color = 2'b11;
		14'h147c: color = 2'b11;
		14'h147d: color = 2'b11;
		14'h147e: color = 2'b11;
		14'h147f: color = 2'b11;
		14'h1480: color = 2'b11;
		14'h1481: color = 2'b11;
		14'h1482: color = 2'b11;
		14'h1483: color = 2'b11;
		14'h1484: color = 2'b11;
		14'h1485: color = 2'b11;
		14'h1486: color = 2'b11;
		14'h1487: color = 2'b11;
		14'h1488: color = 2'b11;
		14'h1489: color = 2'b11;
		14'h148a: color = 2'b11;
		14'h148b: color = 2'b11;
		14'h148c: color = 2'b11;
		14'h148d: color = 2'b11;
		14'h148e: color = 2'b11;
		14'h148f: color = 2'b11;
		14'h1490: color = 2'b11;
		14'h1491: color = 2'b11;
		14'h1492: color = 2'b11;
		14'h1493: color = 2'b11;
		14'h1494: color = 2'b11;
		14'h1495: color = 2'b11;
		14'h1496: color = 2'b11;
		14'h1497: color = 2'b11;
		14'h1498: color = 2'b11;
		14'h1499: color = 2'b11;
		14'h149a: color = 2'b11;
		14'h149b: color = 2'b11;
		14'h149c: color = 2'b11;
		14'h149d: color = 2'b11;
		14'h149e: color = 2'b11;
		14'h149f: color = 2'b11;
		14'h14a0: color = 2'b11;
		14'h14a1: color = 2'b01;
		14'h14a2: color = 2'b01;
		14'h14a3: color = 2'b00;
		14'h14a4: color = 2'b01;
		14'h14a5: color = 2'b00;
		14'h14a6: color = 2'b00;
		14'h14a7: color = 2'b00;
		14'h14a8: color = 2'b00;
		14'h14a9: color = 2'b00;
		14'h14aa: color = 2'b01;
		14'h14ab: color = 2'b01;
		14'h14ac: color = 2'b01;
		14'h14ad: color = 2'b00;
		14'h14ae: color = 2'b01;
		14'h14af: color = 2'b00;
		14'h14b0: color = 2'b01;
		14'h14b1: color = 2'b00;
		14'h14b2: color = 2'b00;
		14'h14b3: color = 2'b00;
		14'h14b4: color = 2'b01;
		14'h14b5: color = 2'b10;
		14'h14b6: color = 2'b11;
		14'h14b7: color = 2'b11;
		14'h14b8: color = 2'b11;
		14'h14b9: color = 2'b11;
		14'h14ba: color = 2'b11;
		14'h14bb: color = 2'b11;
		14'h14bc: color = 2'b11;
		14'h14bd: color = 2'b11;
		14'h14be: color = 2'b11;
		14'h14bf: color = 2'b11;
		14'h14c0: color = 2'b11;
		14'h14c1: color = 2'b11;
		14'h14c2: color = 2'b11;
		14'h14c3: color = 2'b11;
		14'h14c4: color = 2'b10;
		14'h14c5: color = 2'b11;
		14'h14c6: color = 2'b10;
		14'h14c7: color = 2'b10;
		14'h14c8: color = 2'b10;
		14'h14c9: color = 2'b10;
		14'h14ca: color = 2'b10;
		14'h14cb: color = 2'b10;
		14'h14cc: color = 2'b10;
		14'h14cd: color = 2'b10;
		14'h14ce: color = 2'b10;
		14'h14cf: color = 2'b10;
		14'h14d0: color = 2'b10;
		14'h14d1: color = 2'b10;
		14'h14d2: color = 2'b10;
		14'h14d3: color = 2'b11;
		14'h14d4: color = 2'b10;
		14'h14d5: color = 2'b10;
		14'h14d6: color = 2'b10;
		14'h14d7: color = 2'b10;
		14'h14d8: color = 2'b10;
		14'h14d9: color = 2'b10;
		14'h14da: color = 2'b10;
		14'h14db: color = 2'b10;
		14'h14dc: color = 2'b10;
		14'h14dd: color = 2'b10;
		14'h14de: color = 2'b10;
		14'h14df: color = 2'b01;
		14'h14e0: color = 2'b00;
		14'h14e1: color = 2'b00;
		14'h14e2: color = 2'b00;
		14'h14e3: color = 2'b00;
		14'h14e4: color = 2'b00;
		14'h14e5: color = 2'b00;
		14'h14e6: color = 2'b00;
		14'h14e7: color = 2'b00;
		14'h14e8: color = 2'b00;
		14'h14e9: color = 2'b00;
		14'h14ea: color = 2'b01;
		14'h14eb: color = 2'b11;
		14'h14ec: color = 2'b11;
		14'h14ed: color = 2'b11;
		14'h14ee: color = 2'b11;
		14'h14ef: color = 2'b11;
		14'h14f0: color = 2'b11;
		14'h14f1: color = 2'b11;
		14'h14f2: color = 2'b11;
		14'h14f3: color = 2'b11;
		14'h14f4: color = 2'b11;
		14'h14f5: color = 2'b11;
		14'h14f6: color = 2'b11;
		14'h14f7: color = 2'b11;
		14'h14f8: color = 2'b11;
		14'h14f9: color = 2'b11;
		14'h14fa: color = 2'b11;
		14'h14fb: color = 2'b11;
		14'h14fc: color = 2'b11;
		14'h14fd: color = 2'b11;
		14'h14fe: color = 2'b11;
		14'h14ff: color = 2'b11;
		14'h1500: color = 2'b11;
		14'h1501: color = 2'b11;
		14'h1502: color = 2'b11;
		14'h1503: color = 2'b11;
		14'h1504: color = 2'b11;
		14'h1505: color = 2'b11;
		14'h1506: color = 2'b11;
		14'h1507: color = 2'b11;
		14'h1508: color = 2'b11;
		14'h1509: color = 2'b11;
		14'h150a: color = 2'b11;
		14'h150b: color = 2'b11;
		14'h150c: color = 2'b11;
		14'h150d: color = 2'b11;
		14'h150e: color = 2'b11;
		14'h150f: color = 2'b11;
		14'h1510: color = 2'b11;
		14'h1511: color = 2'b11;
		14'h1512: color = 2'b11;
		14'h1513: color = 2'b11;
		14'h1514: color = 2'b11;
		14'h1515: color = 2'b11;
		14'h1516: color = 2'b11;
		14'h1517: color = 2'b11;
		14'h1518: color = 2'b11;
		14'h1519: color = 2'b11;
		14'h151a: color = 2'b11;
		14'h151b: color = 2'b11;
		14'h151c: color = 2'b11;
		14'h151d: color = 2'b11;
		14'h151e: color = 2'b11;
		14'h151f: color = 2'b11;
		14'h1520: color = 2'b10;
		14'h1521: color = 2'b00;
		14'h1522: color = 2'b00;
		14'h1523: color = 2'b00;
		14'h1524: color = 2'b00;
		14'h1525: color = 2'b00;
		14'h1526: color = 2'b00;
		14'h1527: color = 2'b00;
		14'h1528: color = 2'b00;
		14'h1529: color = 2'b01;
		14'h152a: color = 2'b00;
		14'h152b: color = 2'b00;
		14'h152c: color = 2'b00;
		14'h152d: color = 2'b01;
		14'h152e: color = 2'b00;
		14'h152f: color = 2'b00;
		14'h1530: color = 2'b00;
		14'h1531: color = 2'b00;
		14'h1532: color = 2'b01;
		14'h1533: color = 2'b00;
		14'h1534: color = 2'b10;
		14'h1535: color = 2'b11;
		14'h1536: color = 2'b11;
		14'h1537: color = 2'b11;
		14'h1538: color = 2'b11;
		14'h1539: color = 2'b11;
		14'h153a: color = 2'b11;
		14'h153b: color = 2'b11;
		14'h153c: color = 2'b11;
		14'h153d: color = 2'b11;
		14'h153e: color = 2'b11;
		14'h153f: color = 2'b10;
		14'h1540: color = 2'b11;
		14'h1541: color = 2'b11;
		14'h1542: color = 2'b10;
		14'h1543: color = 2'b11;
		14'h1544: color = 2'b11;
		14'h1545: color = 2'b11;
		14'h1546: color = 2'b10;
		14'h1547: color = 2'b11;
		14'h1548: color = 2'b11;
		14'h1549: color = 2'b10;
		14'h154a: color = 2'b10;
		14'h154b: color = 2'b10;
		14'h154c: color = 2'b10;
		14'h154d: color = 2'b10;
		14'h154e: color = 2'b10;
		14'h154f: color = 2'b10;
		14'h1550: color = 2'b10;
		14'h1551: color = 2'b10;
		14'h1552: color = 2'b10;
		14'h1553: color = 2'b10;
		14'h1554: color = 2'b10;
		14'h1555: color = 2'b10;
		14'h1556: color = 2'b10;
		14'h1557: color = 2'b10;
		14'h1558: color = 2'b10;
		14'h1559: color = 2'b10;
		14'h155a: color = 2'b01;
		14'h155b: color = 2'b10;
		14'h155c: color = 2'b01;
		14'h155d: color = 2'b10;
		14'h155e: color = 2'b01;
		14'h155f: color = 2'b10;
		14'h1560: color = 2'b00;
		14'h1561: color = 2'b00;
		14'h1562: color = 2'b00;
		14'h1563: color = 2'b00;
		14'h1564: color = 2'b00;
		14'h1565: color = 2'b00;
		14'h1566: color = 2'b00;
		14'h1567: color = 2'b00;
		14'h1568: color = 2'b00;
		14'h1569: color = 2'b00;
		14'h156a: color = 2'b11;
		14'h156b: color = 2'b11;
		14'h156c: color = 2'b11;
		14'h156d: color = 2'b11;
		14'h156e: color = 2'b11;
		14'h156f: color = 2'b11;
		14'h1570: color = 2'b11;
		14'h1571: color = 2'b11;
		14'h1572: color = 2'b11;
		14'h1573: color = 2'b11;
		14'h1574: color = 2'b11;
		14'h1575: color = 2'b11;
		14'h1576: color = 2'b11;
		14'h1577: color = 2'b11;
		14'h1578: color = 2'b11;
		14'h1579: color = 2'b11;
		14'h157a: color = 2'b11;
		14'h157b: color = 2'b11;
		14'h157c: color = 2'b11;
		14'h157d: color = 2'b11;
		14'h157e: color = 2'b11;
		14'h157f: color = 2'b11;
		14'h1580: color = 2'b11;
		14'h1581: color = 2'b11;
		14'h1582: color = 2'b11;
		14'h1583: color = 2'b11;
		14'h1584: color = 2'b11;
		14'h1585: color = 2'b11;
		14'h1586: color = 2'b11;
		14'h1587: color = 2'b11;
		14'h1588: color = 2'b11;
		14'h1589: color = 2'b11;
		14'h158a: color = 2'b11;
		14'h158b: color = 2'b11;
		14'h158c: color = 2'b11;
		14'h158d: color = 2'b11;
		14'h158e: color = 2'b11;
		14'h158f: color = 2'b11;
		14'h1590: color = 2'b11;
		14'h1591: color = 2'b11;
		14'h1592: color = 2'b11;
		14'h1593: color = 2'b11;
		14'h1594: color = 2'b11;
		14'h1595: color = 2'b11;
		14'h1596: color = 2'b11;
		14'h1597: color = 2'b11;
		14'h1598: color = 2'b11;
		14'h1599: color = 2'b11;
		14'h159a: color = 2'b11;
		14'h159b: color = 2'b11;
		14'h159c: color = 2'b11;
		14'h159d: color = 2'b11;
		14'h159e: color = 2'b11;
		14'h159f: color = 2'b11;
		14'h15a0: color = 2'b10;
		14'h15a1: color = 2'b00;
		14'h15a2: color = 2'b00;
		14'h15a3: color = 2'b00;
		14'h15a4: color = 2'b01;
		14'h15a5: color = 2'b00;
		14'h15a6: color = 2'b00;
		14'h15a7: color = 2'b01;
		14'h15a8: color = 2'b01;
		14'h15a9: color = 2'b00;
		14'h15aa: color = 2'b00;
		14'h15ab: color = 2'b00;
		14'h15ac: color = 2'b00;
		14'h15ad: color = 2'b00;
		14'h15ae: color = 2'b01;
		14'h15af: color = 2'b00;
		14'h15b0: color = 2'b01;
		14'h15b1: color = 2'b00;
		14'h15b2: color = 2'b00;
		14'h15b3: color = 2'b10;
		14'h15b4: color = 2'b11;
		14'h15b5: color = 2'b11;
		14'h15b6: color = 2'b11;
		14'h15b7: color = 2'b11;
		14'h15b8: color = 2'b11;
		14'h15b9: color = 2'b11;
		14'h15ba: color = 2'b11;
		14'h15bb: color = 2'b11;
		14'h15bc: color = 2'b11;
		14'h15bd: color = 2'b11;
		14'h15be: color = 2'b11;
		14'h15bf: color = 2'b11;
		14'h15c0: color = 2'b11;
		14'h15c1: color = 2'b11;
		14'h15c2: color = 2'b11;
		14'h15c3: color = 2'b11;
		14'h15c4: color = 2'b10;
		14'h15c5: color = 2'b11;
		14'h15c6: color = 2'b11;
		14'h15c7: color = 2'b10;
		14'h15c8: color = 2'b10;
		14'h15c9: color = 2'b11;
		14'h15ca: color = 2'b10;
		14'h15cb: color = 2'b10;
		14'h15cc: color = 2'b10;
		14'h15cd: color = 2'b10;
		14'h15ce: color = 2'b10;
		14'h15cf: color = 2'b10;
		14'h15d0: color = 2'b10;
		14'h15d1: color = 2'b11;
		14'h15d2: color = 2'b10;
		14'h15d3: color = 2'b11;
		14'h15d4: color = 2'b10;
		14'h15d5: color = 2'b10;
		14'h15d6: color = 2'b10;
		14'h15d7: color = 2'b10;
		14'h15d8: color = 2'b10;
		14'h15d9: color = 2'b10;
		14'h15da: color = 2'b10;
		14'h15db: color = 2'b10;
		14'h15dc: color = 2'b10;
		14'h15dd: color = 2'b10;
		14'h15de: color = 2'b10;
		14'h15df: color = 2'b01;
		14'h15e0: color = 2'b00;
		14'h15e1: color = 2'b00;
		14'h15e2: color = 2'b00;
		14'h15e3: color = 2'b00;
		14'h15e4: color = 2'b00;
		14'h15e5: color = 2'b00;
		14'h15e6: color = 2'b00;
		14'h15e7: color = 2'b00;
		14'h15e8: color = 2'b00;
		14'h15e9: color = 2'b01;
		14'h15ea: color = 2'b11;
		14'h15eb: color = 2'b11;
		14'h15ec: color = 2'b11;
		14'h15ed: color = 2'b11;
		14'h15ee: color = 2'b11;
		14'h15ef: color = 2'b11;
		14'h15f0: color = 2'b11;
		14'h15f1: color = 2'b11;
		14'h15f2: color = 2'b11;
		14'h15f3: color = 2'b11;
		14'h15f4: color = 2'b11;
		14'h15f5: color = 2'b11;
		14'h15f6: color = 2'b11;
		14'h15f7: color = 2'b11;
		14'h15f8: color = 2'b11;
		14'h15f9: color = 2'b11;
		14'h15fa: color = 2'b11;
		14'h15fb: color = 2'b11;
		14'h15fc: color = 2'b11;
		14'h15fd: color = 2'b11;
		14'h15fe: color = 2'b11;
		14'h15ff: color = 2'b11;
		14'h1600: color = 2'b11;
		14'h1601: color = 2'b11;
		14'h1602: color = 2'b11;
		14'h1603: color = 2'b11;
		14'h1604: color = 2'b11;
		14'h1605: color = 2'b11;
		14'h1606: color = 2'b11;
		14'h1607: color = 2'b11;
		14'h1608: color = 2'b11;
		14'h1609: color = 2'b11;
		14'h160a: color = 2'b11;
		14'h160b: color = 2'b11;
		14'h160c: color = 2'b11;
		14'h160d: color = 2'b11;
		14'h160e: color = 2'b11;
		14'h160f: color = 2'b11;
		14'h1610: color = 2'b11;
		14'h1611: color = 2'b11;
		14'h1612: color = 2'b11;
		14'h1613: color = 2'b11;
		14'h1614: color = 2'b11;
		14'h1615: color = 2'b11;
		14'h1616: color = 2'b11;
		14'h1617: color = 2'b11;
		14'h1618: color = 2'b11;
		14'h1619: color = 2'b11;
		14'h161a: color = 2'b11;
		14'h161b: color = 2'b11;
		14'h161c: color = 2'b11;
		14'h161d: color = 2'b11;
		14'h161e: color = 2'b11;
		14'h161f: color = 2'b11;
		14'h1620: color = 2'b01;
		14'h1621: color = 2'b00;
		14'h1622: color = 2'b00;
		14'h1623: color = 2'b00;
		14'h1624: color = 2'b00;
		14'h1625: color = 2'b01;
		14'h1626: color = 2'b01;
		14'h1627: color = 2'b00;
		14'h1628: color = 2'b00;
		14'h1629: color = 2'b00;
		14'h162a: color = 2'b01;
		14'h162b: color = 2'b00;
		14'h162c: color = 2'b01;
		14'h162d: color = 2'b00;
		14'h162e: color = 2'b00;
		14'h162f: color = 2'b01;
		14'h1630: color = 2'b00;
		14'h1631: color = 2'b00;
		14'h1632: color = 2'b01;
		14'h1633: color = 2'b11;
		14'h1634: color = 2'b11;
		14'h1635: color = 2'b11;
		14'h1636: color = 2'b11;
		14'h1637: color = 2'b11;
		14'h1638: color = 2'b11;
		14'h1639: color = 2'b11;
		14'h163a: color = 2'b11;
		14'h163b: color = 2'b11;
		14'h163c: color = 2'b11;
		14'h163d: color = 2'b11;
		14'h163e: color = 2'b11;
		14'h163f: color = 2'b11;
		14'h1640: color = 2'b10;
		14'h1641: color = 2'b11;
		14'h1642: color = 2'b10;
		14'h1643: color = 2'b11;
		14'h1644: color = 2'b10;
		14'h1645: color = 2'b11;
		14'h1646: color = 2'b10;
		14'h1647: color = 2'b11;
		14'h1648: color = 2'b11;
		14'h1649: color = 2'b10;
		14'h164a: color = 2'b10;
		14'h164b: color = 2'b11;
		14'h164c: color = 2'b10;
		14'h164d: color = 2'b10;
		14'h164e: color = 2'b10;
		14'h164f: color = 2'b10;
		14'h1650: color = 2'b10;
		14'h1651: color = 2'b10;
		14'h1652: color = 2'b10;
		14'h1653: color = 2'b10;
		14'h1654: color = 2'b10;
		14'h1655: color = 2'b10;
		14'h1656: color = 2'b10;
		14'h1657: color = 2'b01;
		14'h1658: color = 2'b01;
		14'h1659: color = 2'b10;
		14'h165a: color = 2'b01;
		14'h165b: color = 2'b10;
		14'h165c: color = 2'b10;
		14'h165d: color = 2'b01;
		14'h165e: color = 2'b10;
		14'h165f: color = 2'b01;
		14'h1660: color = 2'b01;
		14'h1661: color = 2'b00;
		14'h1662: color = 2'b00;
		14'h1663: color = 2'b00;
		14'h1664: color = 2'b00;
		14'h1665: color = 2'b00;
		14'h1666: color = 2'b00;
		14'h1667: color = 2'b00;
		14'h1668: color = 2'b00;
		14'h1669: color = 2'b11;
		14'h166a: color = 2'b11;
		14'h166b: color = 2'b11;
		14'h166c: color = 2'b11;
		14'h166d: color = 2'b11;
		14'h166e: color = 2'b11;
		14'h166f: color = 2'b11;
		14'h1670: color = 2'b11;
		14'h1671: color = 2'b11;
		14'h1672: color = 2'b11;
		14'h1673: color = 2'b11;
		14'h1674: color = 2'b11;
		14'h1675: color = 2'b11;
		14'h1676: color = 2'b11;
		14'h1677: color = 2'b11;
		14'h1678: color = 2'b11;
		14'h1679: color = 2'b11;
		14'h167a: color = 2'b11;
		14'h167b: color = 2'b11;
		14'h167c: color = 2'b11;
		14'h167d: color = 2'b11;
		14'h167e: color = 2'b11;
		14'h167f: color = 2'b11;
		14'h1680: color = 2'b11;
		14'h1681: color = 2'b11;
		14'h1682: color = 2'b11;
		14'h1683: color = 2'b11;
		14'h1684: color = 2'b11;
		14'h1685: color = 2'b11;
		14'h1686: color = 2'b11;
		14'h1687: color = 2'b11;
		14'h1688: color = 2'b11;
		14'h1689: color = 2'b11;
		14'h168a: color = 2'b11;
		14'h168b: color = 2'b11;
		14'h168c: color = 2'b11;
		14'h168d: color = 2'b11;
		14'h168e: color = 2'b11;
		14'h168f: color = 2'b11;
		14'h1690: color = 2'b11;
		14'h1691: color = 2'b11;
		14'h1692: color = 2'b11;
		14'h1693: color = 2'b11;
		14'h1694: color = 2'b11;
		14'h1695: color = 2'b11;
		14'h1696: color = 2'b11;
		14'h1697: color = 2'b11;
		14'h1698: color = 2'b11;
		14'h1699: color = 2'b11;
		14'h169a: color = 2'b11;
		14'h169b: color = 2'b11;
		14'h169c: color = 2'b11;
		14'h169d: color = 2'b11;
		14'h169e: color = 2'b11;
		14'h169f: color = 2'b11;
		14'h16a0: color = 2'b01;
		14'h16a1: color = 2'b00;
		14'h16a2: color = 2'b00;
		14'h16a3: color = 2'b00;
		14'h16a4: color = 2'b01;
		14'h16a5: color = 2'b00;
		14'h16a6: color = 2'b00;
		14'h16a7: color = 2'b00;
		14'h16a8: color = 2'b00;
		14'h16a9: color = 2'b00;
		14'h16aa: color = 2'b00;
		14'h16ab: color = 2'b00;
		14'h16ac: color = 2'b01;
		14'h16ad: color = 2'b00;
		14'h16ae: color = 2'b01;
		14'h16af: color = 2'b00;
		14'h16b0: color = 2'b00;
		14'h16b1: color = 2'b00;
		14'h16b2: color = 2'b10;
		14'h16b3: color = 2'b11;
		14'h16b4: color = 2'b11;
		14'h16b5: color = 2'b11;
		14'h16b6: color = 2'b11;
		14'h16b7: color = 2'b11;
		14'h16b8: color = 2'b11;
		14'h16b9: color = 2'b11;
		14'h16ba: color = 2'b11;
		14'h16bb: color = 2'b11;
		14'h16bc: color = 2'b11;
		14'h16bd: color = 2'b11;
		14'h16be: color = 2'b10;
		14'h16bf: color = 2'b11;
		14'h16c0: color = 2'b10;
		14'h16c1: color = 2'b10;
		14'h16c2: color = 2'b10;
		14'h16c3: color = 2'b10;
		14'h16c4: color = 2'b10;
		14'h16c5: color = 2'b11;
		14'h16c6: color = 2'b10;
		14'h16c7: color = 2'b10;
		14'h16c8: color = 2'b10;
		14'h16c9: color = 2'b11;
		14'h16ca: color = 2'b10;
		14'h16cb: color = 2'b10;
		14'h16cc: color = 2'b10;
		14'h16cd: color = 2'b10;
		14'h16ce: color = 2'b10;
		14'h16cf: color = 2'b10;
		14'h16d0: color = 2'b10;
		14'h16d1: color = 2'b10;
		14'h16d2: color = 2'b10;
		14'h16d3: color = 2'b10;
		14'h16d4: color = 2'b10;
		14'h16d5: color = 2'b01;
		14'h16d6: color = 2'b10;
		14'h16d7: color = 2'b10;
		14'h16d8: color = 2'b10;
		14'h16d9: color = 2'b01;
		14'h16da: color = 2'b10;
		14'h16db: color = 2'b01;
		14'h16dc: color = 2'b01;
		14'h16dd: color = 2'b10;
		14'h16de: color = 2'b01;
		14'h16df: color = 2'b10;
		14'h16e0: color = 2'b00;
		14'h16e1: color = 2'b00;
		14'h16e2: color = 2'b00;
		14'h16e3: color = 2'b00;
		14'h16e4: color = 2'b00;
		14'h16e5: color = 2'b00;
		14'h16e6: color = 2'b10;
		14'h16e7: color = 2'b11;
		14'h16e8: color = 2'b11;
		14'h16e9: color = 2'b11;
		14'h16ea: color = 2'b11;
		14'h16eb: color = 2'b11;
		14'h16ec: color = 2'b11;
		14'h16ed: color = 2'b11;
		14'h16ee: color = 2'b11;
		14'h16ef: color = 2'b11;
		14'h16f0: color = 2'b11;
		14'h16f1: color = 2'b11;
		14'h16f2: color = 2'b11;
		14'h16f3: color = 2'b11;
		14'h16f4: color = 2'b11;
		14'h16f5: color = 2'b11;
		14'h16f6: color = 2'b11;
		14'h16f7: color = 2'b11;
		14'h16f8: color = 2'b11;
		14'h16f9: color = 2'b11;
		14'h16fa: color = 2'b11;
		14'h16fb: color = 2'b11;
		14'h16fc: color = 2'b11;
		14'h16fd: color = 2'b11;
		14'h16fe: color = 2'b11;
		14'h16ff: color = 2'b11;
		14'h1700: color = 2'b11;
		14'h1701: color = 2'b11;
		14'h1702: color = 2'b11;
		14'h1703: color = 2'b11;
		14'h1704: color = 2'b11;
		14'h1705: color = 2'b11;
		14'h1706: color = 2'b11;
		14'h1707: color = 2'b11;
		14'h1708: color = 2'b11;
		14'h1709: color = 2'b11;
		14'h170a: color = 2'b11;
		14'h170b: color = 2'b11;
		14'h170c: color = 2'b11;
		14'h170d: color = 2'b11;
		14'h170e: color = 2'b11;
		14'h170f: color = 2'b11;
		14'h1710: color = 2'b11;
		14'h1711: color = 2'b11;
		14'h1712: color = 2'b11;
		14'h1713: color = 2'b11;
		14'h1714: color = 2'b11;
		14'h1715: color = 2'b11;
		14'h1716: color = 2'b11;
		14'h1717: color = 2'b11;
		14'h1718: color = 2'b11;
		14'h1719: color = 2'b11;
		14'h171a: color = 2'b11;
		14'h171b: color = 2'b11;
		14'h171c: color = 2'b11;
		14'h171d: color = 2'b11;
		14'h171e: color = 2'b11;
		14'h171f: color = 2'b11;
		14'h1720: color = 2'b01;
		14'h1721: color = 2'b00;
		14'h1722: color = 2'b00;
		14'h1723: color = 2'b10;
		14'h1724: color = 2'b01;
		14'h1725: color = 2'b01;
		14'h1726: color = 2'b00;
		14'h1727: color = 2'b01;
		14'h1728: color = 2'b01;
		14'h1729: color = 2'b00;
		14'h172a: color = 2'b00;
		14'h172b: color = 2'b01;
		14'h172c: color = 2'b00;
		14'h172d: color = 2'b01;
		14'h172e: color = 2'b00;
		14'h172f: color = 2'b00;
		14'h1730: color = 2'b01;
		14'h1731: color = 2'b01;
		14'h1732: color = 2'b11;
		14'h1733: color = 2'b11;
		14'h1734: color = 2'b11;
		14'h1735: color = 2'b11;
		14'h1736: color = 2'b11;
		14'h1737: color = 2'b11;
		14'h1738: color = 2'b11;
		14'h1739: color = 2'b11;
		14'h173a: color = 2'b11;
		14'h173b: color = 2'b11;
		14'h173c: color = 2'b11;
		14'h173d: color = 2'b10;
		14'h173e: color = 2'b10;
		14'h173f: color = 2'b10;
		14'h1740: color = 2'b01;
		14'h1741: color = 2'b01;
		14'h1742: color = 2'b01;
		14'h1743: color = 2'b01;
		14'h1744: color = 2'b10;
		14'h1745: color = 2'b01;
		14'h1746: color = 2'b10;
		14'h1747: color = 2'b10;
		14'h1748: color = 2'b10;
		14'h1749: color = 2'b10;
		14'h174a: color = 2'b10;
		14'h174b: color = 2'b10;
		14'h174c: color = 2'b10;
		14'h174d: color = 2'b10;
		14'h174e: color = 2'b10;
		14'h174f: color = 2'b10;
		14'h1750: color = 2'b10;
		14'h1751: color = 2'b10;
		14'h1752: color = 2'b10;
		14'h1753: color = 2'b10;
		14'h1754: color = 2'b01;
		14'h1755: color = 2'b10;
		14'h1756: color = 2'b01;
		14'h1757: color = 2'b10;
		14'h1758: color = 2'b10;
		14'h1759: color = 2'b01;
		14'h175a: color = 2'b01;
		14'h175b: color = 2'b01;
		14'h175c: color = 2'b01;
		14'h175d: color = 2'b01;
		14'h175e: color = 2'b01;
		14'h175f: color = 2'b10;
		14'h1760: color = 2'b00;
		14'h1761: color = 2'b00;
		14'h1762: color = 2'b00;
		14'h1763: color = 2'b00;
		14'h1764: color = 2'b00;
		14'h1765: color = 2'b00;
		14'h1766: color = 2'b11;
		14'h1767: color = 2'b11;
		14'h1768: color = 2'b11;
		14'h1769: color = 2'b11;
		14'h176a: color = 2'b11;
		14'h176b: color = 2'b11;
		14'h176c: color = 2'b11;
		14'h176d: color = 2'b11;
		14'h176e: color = 2'b11;
		14'h176f: color = 2'b11;
		14'h1770: color = 2'b11;
		14'h1771: color = 2'b11;
		14'h1772: color = 2'b11;
		14'h1773: color = 2'b11;
		14'h1774: color = 2'b11;
		14'h1775: color = 2'b11;
		14'h1776: color = 2'b11;
		14'h1777: color = 2'b11;
		14'h1778: color = 2'b11;
		14'h1779: color = 2'b11;
		14'h177a: color = 2'b11;
		14'h177b: color = 2'b11;
		14'h177c: color = 2'b11;
		14'h177d: color = 2'b11;
		14'h177e: color = 2'b11;
		14'h177f: color = 2'b11;
		14'h1780: color = 2'b11;
		14'h1781: color = 2'b11;
		14'h1782: color = 2'b11;
		14'h1783: color = 2'b11;
		14'h1784: color = 2'b11;
		14'h1785: color = 2'b11;
		14'h1786: color = 2'b11;
		14'h1787: color = 2'b11;
		14'h1788: color = 2'b11;
		14'h1789: color = 2'b11;
		14'h178a: color = 2'b11;
		14'h178b: color = 2'b11;
		14'h178c: color = 2'b11;
		14'h178d: color = 2'b11;
		14'h178e: color = 2'b11;
		14'h178f: color = 2'b11;
		14'h1790: color = 2'b11;
		14'h1791: color = 2'b11;
		14'h1792: color = 2'b11;
		14'h1793: color = 2'b11;
		14'h1794: color = 2'b11;
		14'h1795: color = 2'b11;
		14'h1796: color = 2'b11;
		14'h1797: color = 2'b11;
		14'h1798: color = 2'b11;
		14'h1799: color = 2'b11;
		14'h179a: color = 2'b11;
		14'h179b: color = 2'b11;
		14'h179c: color = 2'b11;
		14'h179d: color = 2'b11;
		14'h179e: color = 2'b11;
		14'h179f: color = 2'b11;
		14'h17a0: color = 2'b10;
		14'h17a1: color = 2'b00;
		14'h17a2: color = 2'b10;
		14'h17a3: color = 2'b11;
		14'h17a4: color = 2'b10;
		14'h17a5: color = 2'b01;
		14'h17a6: color = 2'b01;
		14'h17a7: color = 2'b00;
		14'h17a8: color = 2'b00;
		14'h17a9: color = 2'b00;
		14'h17aa: color = 2'b00;
		14'h17ab: color = 2'b00;
		14'h17ac: color = 2'b01;
		14'h17ad: color = 2'b00;
		14'h17ae: color = 2'b00;
		14'h17af: color = 2'b00;
		14'h17b0: color = 2'b01;
		14'h17b1: color = 2'b10;
		14'h17b2: color = 2'b11;
		14'h17b3: color = 2'b11;
		14'h17b4: color = 2'b11;
		14'h17b5: color = 2'b11;
		14'h17b6: color = 2'b11;
		14'h17b7: color = 2'b11;
		14'h17b8: color = 2'b11;
		14'h17b9: color = 2'b11;
		14'h17ba: color = 2'b10;
		14'h17bb: color = 2'b10;
		14'h17bc: color = 2'b01;
		14'h17bd: color = 2'b01;
		14'h17be: color = 2'b01;
		14'h17bf: color = 2'b00;
		14'h17c0: color = 2'b00;
		14'h17c1: color = 2'b00;
		14'h17c2: color = 2'b00;
		14'h17c3: color = 2'b00;
		14'h17c4: color = 2'b00;
		14'h17c5: color = 2'b01;
		14'h17c6: color = 2'b01;
		14'h17c7: color = 2'b01;
		14'h17c8: color = 2'b01;
		14'h17c9: color = 2'b10;
		14'h17ca: color = 2'b01;
		14'h17cb: color = 2'b10;
		14'h17cc: color = 2'b10;
		14'h17cd: color = 2'b10;
		14'h17ce: color = 2'b10;
		14'h17cf: color = 2'b01;
		14'h17d0: color = 2'b01;
		14'h17d1: color = 2'b10;
		14'h17d2: color = 2'b10;
		14'h17d3: color = 2'b01;
		14'h17d4: color = 2'b10;
		14'h17d5: color = 2'b01;
		14'h17d6: color = 2'b01;
		14'h17d7: color = 2'b01;
		14'h17d8: color = 2'b01;
		14'h17d9: color = 2'b01;
		14'h17da: color = 2'b00;
		14'h17db: color = 2'b00;
		14'h17dc: color = 2'b00;
		14'h17dd: color = 2'b00;
		14'h17de: color = 2'b00;
		14'h17df: color = 2'b01;
		14'h17e0: color = 2'b01;
		14'h17e1: color = 2'b00;
		14'h17e2: color = 2'b00;
		14'h17e3: color = 2'b00;
		14'h17e4: color = 2'b00;
		14'h17e5: color = 2'b00;
		14'h17e6: color = 2'b11;
		14'h17e7: color = 2'b11;
		14'h17e8: color = 2'b11;
		14'h17e9: color = 2'b11;
		14'h17ea: color = 2'b11;
		14'h17eb: color = 2'b11;
		14'h17ec: color = 2'b11;
		14'h17ed: color = 2'b11;
		14'h17ee: color = 2'b11;
		14'h17ef: color = 2'b11;
		14'h17f0: color = 2'b11;
		14'h17f1: color = 2'b11;
		14'h17f2: color = 2'b11;
		14'h17f3: color = 2'b11;
		14'h17f4: color = 2'b11;
		14'h17f5: color = 2'b11;
		14'h17f6: color = 2'b11;
		14'h17f7: color = 2'b11;
		14'h17f8: color = 2'b11;
		14'h17f9: color = 2'b11;
		14'h17fa: color = 2'b11;
		14'h17fb: color = 2'b11;
		14'h17fc: color = 2'b11;
		14'h17fd: color = 2'b11;
		14'h17fe: color = 2'b11;
		14'h17ff: color = 2'b11;
		14'h1800: color = 2'b11;
		14'h1801: color = 2'b11;
		14'h1802: color = 2'b11;
		14'h1803: color = 2'b11;
		14'h1804: color = 2'b11;
		14'h1805: color = 2'b11;
		14'h1806: color = 2'b11;
		14'h1807: color = 2'b11;
		14'h1808: color = 2'b11;
		14'h1809: color = 2'b11;
		14'h180a: color = 2'b11;
		14'h180b: color = 2'b11;
		14'h180c: color = 2'b11;
		14'h180d: color = 2'b11;
		14'h180e: color = 2'b11;
		14'h180f: color = 2'b11;
		14'h1810: color = 2'b11;
		14'h1811: color = 2'b11;
		14'h1812: color = 2'b11;
		14'h1813: color = 2'b11;
		14'h1814: color = 2'b11;
		14'h1815: color = 2'b11;
		14'h1816: color = 2'b11;
		14'h1817: color = 2'b11;
		14'h1818: color = 2'b11;
		14'h1819: color = 2'b11;
		14'h181a: color = 2'b11;
		14'h181b: color = 2'b11;
		14'h181c: color = 2'b11;
		14'h181d: color = 2'b11;
		14'h181e: color = 2'b11;
		14'h181f: color = 2'b11;
		14'h1820: color = 2'b10;
		14'h1821: color = 2'b10;
		14'h1822: color = 2'b10;
		14'h1823: color = 2'b10;
		14'h1824: color = 2'b10;
		14'h1825: color = 2'b11;
		14'h1826: color = 2'b11;
		14'h1827: color = 2'b10;
		14'h1828: color = 2'b10;
		14'h1829: color = 2'b01;
		14'h182a: color = 2'b00;
		14'h182b: color = 2'b00;
		14'h182c: color = 2'b00;
		14'h182d: color = 2'b00;
		14'h182e: color = 2'b00;
		14'h182f: color = 2'b00;
		14'h1830: color = 2'b01;
		14'h1831: color = 2'b11;
		14'h1832: color = 2'b11;
		14'h1833: color = 2'b11;
		14'h1834: color = 2'b11;
		14'h1835: color = 2'b11;
		14'h1836: color = 2'b11;
		14'h1837: color = 2'b11;
		14'h1838: color = 2'b11;
		14'h1839: color = 2'b11;
		14'h183a: color = 2'b10;
		14'h183b: color = 2'b10;
		14'h183c: color = 2'b10;
		14'h183d: color = 2'b01;
		14'h183e: color = 2'b01;
		14'h183f: color = 2'b01;
		14'h1840: color = 2'b01;
		14'h1841: color = 2'b00;
		14'h1842: color = 2'b00;
		14'h1843: color = 2'b00;
		14'h1844: color = 2'b00;
		14'h1845: color = 2'b00;
		14'h1846: color = 2'b00;
		14'h1847: color = 2'b00;
		14'h1848: color = 2'b00;
		14'h1849: color = 2'b00;
		14'h184a: color = 2'b01;
		14'h184b: color = 2'b01;
		14'h184c: color = 2'b01;
		14'h184d: color = 2'b01;
		14'h184e: color = 2'b10;
		14'h184f: color = 2'b01;
		14'h1850: color = 2'b01;
		14'h1851: color = 2'b01;
		14'h1852: color = 2'b01;
		14'h1853: color = 2'b01;
		14'h1854: color = 2'b01;
		14'h1855: color = 2'b00;
		14'h1856: color = 2'b00;
		14'h1857: color = 2'b00;
		14'h1858: color = 2'b00;
		14'h1859: color = 2'b00;
		14'h185a: color = 2'b00;
		14'h185b: color = 2'b00;
		14'h185c: color = 2'b00;
		14'h185d: color = 2'b00;
		14'h185e: color = 2'b00;
		14'h185f: color = 2'b00;
		14'h1860: color = 2'b01;
		14'h1861: color = 2'b00;
		14'h1862: color = 2'b00;
		14'h1863: color = 2'b00;
		14'h1864: color = 2'b00;
		14'h1865: color = 2'b00;
		14'h1866: color = 2'b11;
		14'h1867: color = 2'b11;
		14'h1868: color = 2'b11;
		14'h1869: color = 2'b11;
		14'h186a: color = 2'b11;
		14'h186b: color = 2'b11;
		14'h186c: color = 2'b11;
		14'h186d: color = 2'b11;
		14'h186e: color = 2'b11;
		14'h186f: color = 2'b11;
		14'h1870: color = 2'b11;
		14'h1871: color = 2'b11;
		14'h1872: color = 2'b11;
		14'h1873: color = 2'b11;
		14'h1874: color = 2'b11;
		14'h1875: color = 2'b11;
		14'h1876: color = 2'b11;
		14'h1877: color = 2'b11;
		14'h1878: color = 2'b11;
		14'h1879: color = 2'b11;
		14'h187a: color = 2'b11;
		14'h187b: color = 2'b11;
		14'h187c: color = 2'b11;
		14'h187d: color = 2'b11;
		14'h187e: color = 2'b11;
		14'h187f: color = 2'b11;
		14'h1880: color = 2'b11;
		14'h1881: color = 2'b11;
		14'h1882: color = 2'b11;
		14'h1883: color = 2'b11;
		14'h1884: color = 2'b11;
		14'h1885: color = 2'b11;
		14'h1886: color = 2'b11;
		14'h1887: color = 2'b11;
		14'h1888: color = 2'b11;
		14'h1889: color = 2'b11;
		14'h188a: color = 2'b11;
		14'h188b: color = 2'b11;
		14'h188c: color = 2'b11;
		14'h188d: color = 2'b11;
		14'h188e: color = 2'b11;
		14'h188f: color = 2'b11;
		14'h1890: color = 2'b11;
		14'h1891: color = 2'b11;
		14'h1892: color = 2'b11;
		14'h1893: color = 2'b11;
		14'h1894: color = 2'b11;
		14'h1895: color = 2'b11;
		14'h1896: color = 2'b11;
		14'h1897: color = 2'b11;
		14'h1898: color = 2'b11;
		14'h1899: color = 2'b11;
		14'h189a: color = 2'b11;
		14'h189b: color = 2'b11;
		14'h189c: color = 2'b11;
		14'h189d: color = 2'b11;
		14'h189e: color = 2'b11;
		14'h189f: color = 2'b11;
		14'h18a0: color = 2'b11;
		14'h18a1: color = 2'b11;
		14'h18a2: color = 2'b01;
		14'h18a3: color = 2'b01;
		14'h18a4: color = 2'b10;
		14'h18a5: color = 2'b10;
		14'h18a6: color = 2'b10;
		14'h18a7: color = 2'b10;
		14'h18a8: color = 2'b10;
		14'h18a9: color = 2'b01;
		14'h18aa: color = 2'b01;
		14'h18ab: color = 2'b00;
		14'h18ac: color = 2'b00;
		14'h18ad: color = 2'b00;
		14'h18ae: color = 2'b01;
		14'h18af: color = 2'b01;
		14'h18b0: color = 2'b01;
		14'h18b1: color = 2'b10;
		14'h18b2: color = 2'b10;
		14'h18b3: color = 2'b11;
		14'h18b4: color = 2'b11;
		14'h18b5: color = 2'b11;
		14'h18b6: color = 2'b11;
		14'h18b7: color = 2'b11;
		14'h18b8: color = 2'b11;
		14'h18b9: color = 2'b10;
		14'h18ba: color = 2'b11;
		14'h18bb: color = 2'b10;
		14'h18bc: color = 2'b10;
		14'h18bd: color = 2'b10;
		14'h18be: color = 2'b10;
		14'h18bf: color = 2'b01;
		14'h18c0: color = 2'b01;
		14'h18c1: color = 2'b01;
		14'h18c2: color = 2'b01;
		14'h18c3: color = 2'b01;
		14'h18c4: color = 2'b01;
		14'h18c5: color = 2'b01;
		14'h18c6: color = 2'b00;
		14'h18c7: color = 2'b01;
		14'h18c8: color = 2'b01;
		14'h18c9: color = 2'b00;
		14'h18ca: color = 2'b00;
		14'h18cb: color = 2'b00;
		14'h18cc: color = 2'b01;
		14'h18cd: color = 2'b01;
		14'h18ce: color = 2'b10;
		14'h18cf: color = 2'b01;
		14'h18d0: color = 2'b01;
		14'h18d1: color = 2'b01;
		14'h18d2: color = 2'b00;
		14'h18d3: color = 2'b00;
		14'h18d4: color = 2'b00;
		14'h18d5: color = 2'b00;
		14'h18d6: color = 2'b00;
		14'h18d7: color = 2'b00;
		14'h18d8: color = 2'b00;
		14'h18d9: color = 2'b00;
		14'h18da: color = 2'b00;
		14'h18db: color = 2'b00;
		14'h18dc: color = 2'b00;
		14'h18dd: color = 2'b01;
		14'h18de: color = 2'b00;
		14'h18df: color = 2'b00;
		14'h18e0: color = 2'b01;
		14'h18e1: color = 2'b00;
		14'h18e2: color = 2'b00;
		14'h18e3: color = 2'b00;
		14'h18e4: color = 2'b00;
		14'h18e5: color = 2'b01;
		14'h18e6: color = 2'b11;
		14'h18e7: color = 2'b11;
		14'h18e8: color = 2'b11;
		14'h18e9: color = 2'b11;
		14'h18ea: color = 2'b11;
		14'h18eb: color = 2'b11;
		14'h18ec: color = 2'b11;
		14'h18ed: color = 2'b11;
		14'h18ee: color = 2'b11;
		14'h18ef: color = 2'b11;
		14'h18f0: color = 2'b11;
		14'h18f1: color = 2'b11;
		14'h18f2: color = 2'b11;
		14'h18f3: color = 2'b11;
		14'h18f4: color = 2'b11;
		14'h18f5: color = 2'b11;
		14'h18f6: color = 2'b11;
		14'h18f7: color = 2'b11;
		14'h18f8: color = 2'b11;
		14'h18f9: color = 2'b11;
		14'h18fa: color = 2'b11;
		14'h18fb: color = 2'b11;
		14'h18fc: color = 2'b11;
		14'h18fd: color = 2'b11;
		14'h18fe: color = 2'b11;
		14'h18ff: color = 2'b11;
		14'h1900: color = 2'b11;
		14'h1901: color = 2'b11;
		14'h1902: color = 2'b11;
		14'h1903: color = 2'b11;
		14'h1904: color = 2'b11;
		14'h1905: color = 2'b11;
		14'h1906: color = 2'b11;
		14'h1907: color = 2'b11;
		14'h1908: color = 2'b11;
		14'h1909: color = 2'b11;
		14'h190a: color = 2'b11;
		14'h190b: color = 2'b11;
		14'h190c: color = 2'b11;
		14'h190d: color = 2'b11;
		14'h190e: color = 2'b11;
		14'h190f: color = 2'b11;
		14'h1910: color = 2'b11;
		14'h1911: color = 2'b11;
		14'h1912: color = 2'b11;
		14'h1913: color = 2'b11;
		14'h1914: color = 2'b11;
		14'h1915: color = 2'b11;
		14'h1916: color = 2'b11;
		14'h1917: color = 2'b11;
		14'h1918: color = 2'b11;
		14'h1919: color = 2'b11;
		14'h191a: color = 2'b11;
		14'h191b: color = 2'b11;
		14'h191c: color = 2'b11;
		14'h191d: color = 2'b11;
		14'h191e: color = 2'b11;
		14'h191f: color = 2'b11;
		14'h1920: color = 2'b10;
		14'h1921: color = 2'b11;
		14'h1922: color = 2'b10;
		14'h1923: color = 2'b10;
		14'h1924: color = 2'b11;
		14'h1925: color = 2'b11;
		14'h1926: color = 2'b10;
		14'h1927: color = 2'b10;
		14'h1928: color = 2'b10;
		14'h1929: color = 2'b10;
		14'h192a: color = 2'b01;
		14'h192b: color = 2'b00;
		14'h192c: color = 2'b01;
		14'h192d: color = 2'b00;
		14'h192e: color = 2'b00;
		14'h192f: color = 2'b01;
		14'h1930: color = 2'b10;
		14'h1931: color = 2'b10;
		14'h1932: color = 2'b10;
		14'h1933: color = 2'b10;
		14'h1934: color = 2'b10;
		14'h1935: color = 2'b11;
		14'h1936: color = 2'b11;
		14'h1937: color = 2'b10;
		14'h1938: color = 2'b10;
		14'h1939: color = 2'b10;
		14'h193a: color = 2'b10;
		14'h193b: color = 2'b11;
		14'h193c: color = 2'b10;
		14'h193d: color = 2'b10;
		14'h193e: color = 2'b01;
		14'h193f: color = 2'b01;
		14'h1940: color = 2'b01;
		14'h1941: color = 2'b01;
		14'h1942: color = 2'b01;
		14'h1943: color = 2'b01;
		14'h1944: color = 2'b01;
		14'h1945: color = 2'b01;
		14'h1946: color = 2'b01;
		14'h1947: color = 2'b01;
		14'h1948: color = 2'b01;
		14'h1949: color = 2'b01;
		14'h194a: color = 2'b01;
		14'h194b: color = 2'b10;
		14'h194c: color = 2'b01;
		14'h194d: color = 2'b10;
		14'h194e: color = 2'b01;
		14'h194f: color = 2'b01;
		14'h1950: color = 2'b01;
		14'h1951: color = 2'b00;
		14'h1952: color = 2'b00;
		14'h1953: color = 2'b00;
		14'h1954: color = 2'b00;
		14'h1955: color = 2'b01;
		14'h1956: color = 2'b00;
		14'h1957: color = 2'b01;
		14'h1958: color = 2'b01;
		14'h1959: color = 2'b01;
		14'h195a: color = 2'b01;
		14'h195b: color = 2'b01;
		14'h195c: color = 2'b01;
		14'h195d: color = 2'b01;
		14'h195e: color = 2'b01;
		14'h195f: color = 2'b01;
		14'h1960: color = 2'b01;
		14'h1961: color = 2'b00;
		14'h1962: color = 2'b00;
		14'h1963: color = 2'b00;
		14'h1964: color = 2'b00;
		14'h1965: color = 2'b11;
		14'h1966: color = 2'b11;
		14'h1967: color = 2'b11;
		14'h1968: color = 2'b11;
		14'h1969: color = 2'b11;
		14'h196a: color = 2'b11;
		14'h196b: color = 2'b11;
		14'h196c: color = 2'b11;
		14'h196d: color = 2'b11;
		14'h196e: color = 2'b11;
		14'h196f: color = 2'b11;
		14'h1970: color = 2'b11;
		14'h1971: color = 2'b11;
		14'h1972: color = 2'b11;
		14'h1973: color = 2'b11;
		14'h1974: color = 2'b11;
		14'h1975: color = 2'b11;
		14'h1976: color = 2'b11;
		14'h1977: color = 2'b11;
		14'h1978: color = 2'b11;
		14'h1979: color = 2'b11;
		14'h197a: color = 2'b11;
		14'h197b: color = 2'b11;
		14'h197c: color = 2'b11;
		14'h197d: color = 2'b11;
		14'h197e: color = 2'b11;
		14'h197f: color = 2'b11;
		14'h1980: color = 2'b11;
		14'h1981: color = 2'b11;
		14'h1982: color = 2'b11;
		14'h1983: color = 2'b11;
		14'h1984: color = 2'b11;
		14'h1985: color = 2'b11;
		14'h1986: color = 2'b11;
		14'h1987: color = 2'b11;
		14'h1988: color = 2'b11;
		14'h1989: color = 2'b11;
		14'h198a: color = 2'b11;
		14'h198b: color = 2'b11;
		14'h198c: color = 2'b11;
		14'h198d: color = 2'b11;
		14'h198e: color = 2'b11;
		14'h198f: color = 2'b11;
		14'h1990: color = 2'b11;
		14'h1991: color = 2'b11;
		14'h1992: color = 2'b11;
		14'h1993: color = 2'b11;
		14'h1994: color = 2'b11;
		14'h1995: color = 2'b11;
		14'h1996: color = 2'b11;
		14'h1997: color = 2'b11;
		14'h1998: color = 2'b11;
		14'h1999: color = 2'b11;
		14'h199a: color = 2'b11;
		14'h199b: color = 2'b11;
		14'h199c: color = 2'b11;
		14'h199d: color = 2'b11;
		14'h199e: color = 2'b11;
		14'h199f: color = 2'b11;
		14'h19a0: color = 2'b11;
		14'h19a1: color = 2'b11;
		14'h19a2: color = 2'b10;
		14'h19a3: color = 2'b10;
		14'h19a4: color = 2'b11;
		14'h19a5: color = 2'b11;
		14'h19a6: color = 2'b11;
		14'h19a7: color = 2'b10;
		14'h19a8: color = 2'b10;
		14'h19a9: color = 2'b10;
		14'h19aa: color = 2'b01;
		14'h19ab: color = 2'b00;
		14'h19ac: color = 2'b00;
		14'h19ad: color = 2'b01;
		14'h19ae: color = 2'b00;
		14'h19af: color = 2'b01;
		14'h19b0: color = 2'b11;
		14'h19b1: color = 2'b11;
		14'h19b2: color = 2'b11;
		14'h19b3: color = 2'b10;
		14'h19b4: color = 2'b10;
		14'h19b5: color = 2'b10;
		14'h19b6: color = 2'b10;
		14'h19b7: color = 2'b10;
		14'h19b8: color = 2'b10;
		14'h19b9: color = 2'b10;
		14'h19ba: color = 2'b10;
		14'h19bb: color = 2'b10;
		14'h19bc: color = 2'b01;
		14'h19bd: color = 2'b01;
		14'h19be: color = 2'b01;
		14'h19bf: color = 2'b01;
		14'h19c0: color = 2'b01;
		14'h19c1: color = 2'b00;
		14'h19c2: color = 2'b00;
		14'h19c3: color = 2'b00;
		14'h19c4: color = 2'b00;
		14'h19c5: color = 2'b00;
		14'h19c6: color = 2'b01;
		14'h19c7: color = 2'b01;
		14'h19c8: color = 2'b01;
		14'h19c9: color = 2'b01;
		14'h19ca: color = 2'b10;
		14'h19cb: color = 2'b10;
		14'h19cc: color = 2'b10;
		14'h19cd: color = 2'b10;
		14'h19ce: color = 2'b01;
		14'h19cf: color = 2'b10;
		14'h19d0: color = 2'b01;
		14'h19d1: color = 2'b01;
		14'h19d2: color = 2'b00;
		14'h19d3: color = 2'b00;
		14'h19d4: color = 2'b00;
		14'h19d5: color = 2'b00;
		14'h19d6: color = 2'b00;
		14'h19d7: color = 2'b00;
		14'h19d8: color = 2'b00;
		14'h19d9: color = 2'b00;
		14'h19da: color = 2'b00;
		14'h19db: color = 2'b00;
		14'h19dc: color = 2'b00;
		14'h19dd: color = 2'b01;
		14'h19de: color = 2'b01;
		14'h19df: color = 2'b01;
		14'h19e0: color = 2'b00;
		14'h19e1: color = 2'b00;
		14'h19e2: color = 2'b00;
		14'h19e3: color = 2'b00;
		14'h19e4: color = 2'b00;
		14'h19e5: color = 2'b11;
		14'h19e6: color = 2'b11;
		14'h19e7: color = 2'b11;
		14'h19e8: color = 2'b11;
		14'h19e9: color = 2'b11;
		14'h19ea: color = 2'b11;
		14'h19eb: color = 2'b11;
		14'h19ec: color = 2'b11;
		14'h19ed: color = 2'b11;
		14'h19ee: color = 2'b11;
		14'h19ef: color = 2'b11;
		14'h19f0: color = 2'b11;
		14'h19f1: color = 2'b11;
		14'h19f2: color = 2'b11;
		14'h19f3: color = 2'b11;
		14'h19f4: color = 2'b11;
		14'h19f5: color = 2'b11;
		14'h19f6: color = 2'b11;
		14'h19f7: color = 2'b11;
		14'h19f8: color = 2'b11;
		14'h19f9: color = 2'b11;
		14'h19fa: color = 2'b11;
		14'h19fb: color = 2'b11;
		14'h19fc: color = 2'b11;
		14'h19fd: color = 2'b11;
		14'h19fe: color = 2'b11;
		14'h19ff: color = 2'b11;
		14'h1a00: color = 2'b11;
		14'h1a01: color = 2'b11;
		14'h1a02: color = 2'b11;
		14'h1a03: color = 2'b11;
		14'h1a04: color = 2'b11;
		14'h1a05: color = 2'b11;
		14'h1a06: color = 2'b11;
		14'h1a07: color = 2'b11;
		14'h1a08: color = 2'b11;
		14'h1a09: color = 2'b11;
		14'h1a0a: color = 2'b11;
		14'h1a0b: color = 2'b11;
		14'h1a0c: color = 2'b11;
		14'h1a0d: color = 2'b11;
		14'h1a0e: color = 2'b11;
		14'h1a0f: color = 2'b11;
		14'h1a10: color = 2'b11;
		14'h1a11: color = 2'b11;
		14'h1a12: color = 2'b11;
		14'h1a13: color = 2'b11;
		14'h1a14: color = 2'b11;
		14'h1a15: color = 2'b11;
		14'h1a16: color = 2'b11;
		14'h1a17: color = 2'b11;
		14'h1a18: color = 2'b11;
		14'h1a19: color = 2'b11;
		14'h1a1a: color = 2'b11;
		14'h1a1b: color = 2'b11;
		14'h1a1c: color = 2'b11;
		14'h1a1d: color = 2'b11;
		14'h1a1e: color = 2'b11;
		14'h1a1f: color = 2'b11;
		14'h1a20: color = 2'b11;
		14'h1a21: color = 2'b11;
		14'h1a22: color = 2'b10;
		14'h1a23: color = 2'b10;
		14'h1a24: color = 2'b11;
		14'h1a25: color = 2'b11;
		14'h1a26: color = 2'b10;
		14'h1a27: color = 2'b10;
		14'h1a28: color = 2'b10;
		14'h1a29: color = 2'b01;
		14'h1a2a: color = 2'b01;
		14'h1a2b: color = 2'b01;
		14'h1a2c: color = 2'b01;
		14'h1a2d: color = 2'b00;
		14'h1a2e: color = 2'b00;
		14'h1a2f: color = 2'b01;
		14'h1a30: color = 2'b10;
		14'h1a31: color = 2'b11;
		14'h1a32: color = 2'b11;
		14'h1a33: color = 2'b11;
		14'h1a34: color = 2'b11;
		14'h1a35: color = 2'b01;
		14'h1a36: color = 2'b10;
		14'h1a37: color = 2'b10;
		14'h1a38: color = 2'b10;
		14'h1a39: color = 2'b10;
		14'h1a3a: color = 2'b10;
		14'h1a3b: color = 2'b10;
		14'h1a3c: color = 2'b01;
		14'h1a3d: color = 2'b10;
		14'h1a3e: color = 2'b01;
		14'h1a3f: color = 2'b10;
		14'h1a40: color = 2'b01;
		14'h1a41: color = 2'b00;
		14'h1a42: color = 2'b00;
		14'h1a43: color = 2'b01;
		14'h1a44: color = 2'b01;
		14'h1a45: color = 2'b01;
		14'h1a46: color = 2'b00;
		14'h1a47: color = 2'b00;
		14'h1a48: color = 2'b00;
		14'h1a49: color = 2'b01;
		14'h1a4a: color = 2'b10;
		14'h1a4b: color = 2'b10;
		14'h1a4c: color = 2'b01;
		14'h1a4d: color = 2'b01;
		14'h1a4e: color = 2'b10;
		14'h1a4f: color = 2'b01;
		14'h1a50: color = 2'b01;
		14'h1a51: color = 2'b01;
		14'h1a52: color = 2'b00;
		14'h1a53: color = 2'b00;
		14'h1a54: color = 2'b00;
		14'h1a55: color = 2'b00;
		14'h1a56: color = 2'b00;
		14'h1a57: color = 2'b00;
		14'h1a58: color = 2'b00;
		14'h1a59: color = 2'b00;
		14'h1a5a: color = 2'b00;
		14'h1a5b: color = 2'b00;
		14'h1a5c: color = 2'b00;
		14'h1a5d: color = 2'b01;
		14'h1a5e: color = 2'b01;
		14'h1a5f: color = 2'b00;
		14'h1a60: color = 2'b00;
		14'h1a61: color = 2'b00;
		14'h1a62: color = 2'b00;
		14'h1a63: color = 2'b00;
		14'h1a64: color = 2'b11;
		14'h1a65: color = 2'b11;
		14'h1a66: color = 2'b11;
		14'h1a67: color = 2'b11;
		14'h1a68: color = 2'b11;
		14'h1a69: color = 2'b11;
		14'h1a6a: color = 2'b11;
		14'h1a6b: color = 2'b11;
		14'h1a6c: color = 2'b11;
		14'h1a6d: color = 2'b11;
		14'h1a6e: color = 2'b11;
		14'h1a6f: color = 2'b11;
		14'h1a70: color = 2'b11;
		14'h1a71: color = 2'b11;
		14'h1a72: color = 2'b11;
		14'h1a73: color = 2'b11;
		14'h1a74: color = 2'b11;
		14'h1a75: color = 2'b11;
		14'h1a76: color = 2'b11;
		14'h1a77: color = 2'b11;
		14'h1a78: color = 2'b11;
		14'h1a79: color = 2'b11;
		14'h1a7a: color = 2'b11;
		14'h1a7b: color = 2'b11;
		14'h1a7c: color = 2'b11;
		14'h1a7d: color = 2'b11;
		14'h1a7e: color = 2'b11;
		14'h1a7f: color = 2'b11;
		14'h1a80: color = 2'b11;
		14'h1a81: color = 2'b11;
		14'h1a82: color = 2'b11;
		14'h1a83: color = 2'b11;
		14'h1a84: color = 2'b11;
		14'h1a85: color = 2'b11;
		14'h1a86: color = 2'b11;
		14'h1a87: color = 2'b11;
		14'h1a88: color = 2'b11;
		14'h1a89: color = 2'b11;
		14'h1a8a: color = 2'b11;
		14'h1a8b: color = 2'b11;
		14'h1a8c: color = 2'b11;
		14'h1a8d: color = 2'b11;
		14'h1a8e: color = 2'b11;
		14'h1a8f: color = 2'b11;
		14'h1a90: color = 2'b11;
		14'h1a91: color = 2'b11;
		14'h1a92: color = 2'b11;
		14'h1a93: color = 2'b11;
		14'h1a94: color = 2'b11;
		14'h1a95: color = 2'b11;
		14'h1a96: color = 2'b11;
		14'h1a97: color = 2'b11;
		14'h1a98: color = 2'b11;
		14'h1a99: color = 2'b11;
		14'h1a9a: color = 2'b11;
		14'h1a9b: color = 2'b11;
		14'h1a9c: color = 2'b11;
		14'h1a9d: color = 2'b11;
		14'h1a9e: color = 2'b11;
		14'h1a9f: color = 2'b11;
		14'h1aa0: color = 2'b11;
		14'h1aa1: color = 2'b11;
		14'h1aa2: color = 2'b01;
		14'h1aa3: color = 2'b10;
		14'h1aa4: color = 2'b11;
		14'h1aa5: color = 2'b11;
		14'h1aa6: color = 2'b10;
		14'h1aa7: color = 2'b10;
		14'h1aa8: color = 2'b10;
		14'h1aa9: color = 2'b01;
		14'h1aaa: color = 2'b01;
		14'h1aab: color = 2'b00;
		14'h1aac: color = 2'b01;
		14'h1aad: color = 2'b00;
		14'h1aae: color = 2'b01;
		14'h1aaf: color = 2'b01;
		14'h1ab0: color = 2'b11;
		14'h1ab1: color = 2'b11;
		14'h1ab2: color = 2'b11;
		14'h1ab3: color = 2'b11;
		14'h1ab4: color = 2'b11;
		14'h1ab5: color = 2'b11;
		14'h1ab6: color = 2'b11;
		14'h1ab7: color = 2'b10;
		14'h1ab8: color = 2'b10;
		14'h1ab9: color = 2'b10;
		14'h1aba: color = 2'b01;
		14'h1abb: color = 2'b10;
		14'h1abc: color = 2'b10;
		14'h1abd: color = 2'b11;
		14'h1abe: color = 2'b10;
		14'h1abf: color = 2'b10;
		14'h1ac0: color = 2'b01;
		14'h1ac1: color = 2'b00;
		14'h1ac2: color = 2'b10;
		14'h1ac3: color = 2'b01;
		14'h1ac4: color = 2'b10;
		14'h1ac5: color = 2'b01;
		14'h1ac6: color = 2'b01;
		14'h1ac7: color = 2'b01;
		14'h1ac8: color = 2'b01;
		14'h1ac9: color = 2'b10;
		14'h1aca: color = 2'b10;
		14'h1acb: color = 2'b01;
		14'h1acc: color = 2'b01;
		14'h1acd: color = 2'b01;
		14'h1ace: color = 2'b10;
		14'h1acf: color = 2'b01;
		14'h1ad0: color = 2'b01;
		14'h1ad1: color = 2'b01;
		14'h1ad2: color = 2'b01;
		14'h1ad3: color = 2'b00;
		14'h1ad4: color = 2'b00;
		14'h1ad5: color = 2'b00;
		14'h1ad6: color = 2'b00;
		14'h1ad7: color = 2'b00;
		14'h1ad8: color = 2'b00;
		14'h1ad9: color = 2'b01;
		14'h1ada: color = 2'b01;
		14'h1adb: color = 2'b01;
		14'h1adc: color = 2'b00;
		14'h1add: color = 2'b01;
		14'h1ade: color = 2'b00;
		14'h1adf: color = 2'b01;
		14'h1ae0: color = 2'b00;
		14'h1ae1: color = 2'b01;
		14'h1ae2: color = 2'b00;
		14'h1ae3: color = 2'b10;
		14'h1ae4: color = 2'b11;
		14'h1ae5: color = 2'b11;
		14'h1ae6: color = 2'b11;
		14'h1ae7: color = 2'b11;
		14'h1ae8: color = 2'b11;
		14'h1ae9: color = 2'b11;
		14'h1aea: color = 2'b11;
		14'h1aeb: color = 2'b11;
		14'h1aec: color = 2'b11;
		14'h1aed: color = 2'b11;
		14'h1aee: color = 2'b11;
		14'h1aef: color = 2'b11;
		14'h1af0: color = 2'b11;
		14'h1af1: color = 2'b11;
		14'h1af2: color = 2'b11;
		14'h1af3: color = 2'b11;
		14'h1af4: color = 2'b11;
		14'h1af5: color = 2'b11;
		14'h1af6: color = 2'b11;
		14'h1af7: color = 2'b11;
		14'h1af8: color = 2'b11;
		14'h1af9: color = 2'b11;
		14'h1afa: color = 2'b11;
		14'h1afb: color = 2'b11;
		14'h1afc: color = 2'b11;
		14'h1afd: color = 2'b11;
		14'h1afe: color = 2'b11;
		14'h1aff: color = 2'b11;
		14'h1b00: color = 2'b11;
		14'h1b01: color = 2'b11;
		14'h1b02: color = 2'b11;
		14'h1b03: color = 2'b11;
		14'h1b04: color = 2'b11;
		14'h1b05: color = 2'b11;
		14'h1b06: color = 2'b11;
		14'h1b07: color = 2'b11;
		14'h1b08: color = 2'b11;
		14'h1b09: color = 2'b11;
		14'h1b0a: color = 2'b11;
		14'h1b0b: color = 2'b11;
		14'h1b0c: color = 2'b11;
		14'h1b0d: color = 2'b11;
		14'h1b0e: color = 2'b11;
		14'h1b0f: color = 2'b11;
		14'h1b10: color = 2'b11;
		14'h1b11: color = 2'b11;
		14'h1b12: color = 2'b11;
		14'h1b13: color = 2'b11;
		14'h1b14: color = 2'b11;
		14'h1b15: color = 2'b11;
		14'h1b16: color = 2'b11;
		14'h1b17: color = 2'b11;
		14'h1b18: color = 2'b11;
		14'h1b19: color = 2'b11;
		14'h1b1a: color = 2'b11;
		14'h1b1b: color = 2'b11;
		14'h1b1c: color = 2'b11;
		14'h1b1d: color = 2'b11;
		14'h1b1e: color = 2'b11;
		14'h1b1f: color = 2'b11;
		14'h1b20: color = 2'b11;
		14'h1b21: color = 2'b11;
		14'h1b22: color = 2'b10;
		14'h1b23: color = 2'b01;
		14'h1b24: color = 2'b10;
		14'h1b25: color = 2'b11;
		14'h1b26: color = 2'b10;
		14'h1b27: color = 2'b10;
		14'h1b28: color = 2'b10;
		14'h1b29: color = 2'b01;
		14'h1b2a: color = 2'b01;
		14'h1b2b: color = 2'b00;
		14'h1b2c: color = 2'b00;
		14'h1b2d: color = 2'b01;
		14'h1b2e: color = 2'b00;
		14'h1b2f: color = 2'b10;
		14'h1b30: color = 2'b11;
		14'h1b31: color = 2'b11;
		14'h1b32: color = 2'b11;
		14'h1b33: color = 2'b11;
		14'h1b34: color = 2'b11;
		14'h1b35: color = 2'b11;
		14'h1b36: color = 2'b11;
		14'h1b37: color = 2'b11;
		14'h1b38: color = 2'b11;
		14'h1b39: color = 2'b10;
		14'h1b3a: color = 2'b10;
		14'h1b3b: color = 2'b10;
		14'h1b3c: color = 2'b11;
		14'h1b3d: color = 2'b10;
		14'h1b3e: color = 2'b10;
		14'h1b3f: color = 2'b11;
		14'h1b40: color = 2'b10;
		14'h1b41: color = 2'b10;
		14'h1b42: color = 2'b01;
		14'h1b43: color = 2'b01;
		14'h1b44: color = 2'b10;
		14'h1b45: color = 2'b01;
		14'h1b46: color = 2'b10;
		14'h1b47: color = 2'b01;
		14'h1b48: color = 2'b01;
		14'h1b49: color = 2'b01;
		14'h1b4a: color = 2'b01;
		14'h1b4b: color = 2'b01;
		14'h1b4c: color = 2'b01;
		14'h1b4d: color = 2'b11;
		14'h1b4e: color = 2'b10;
		14'h1b4f: color = 2'b10;
		14'h1b50: color = 2'b01;
		14'h1b51: color = 2'b00;
		14'h1b52: color = 2'b01;
		14'h1b53: color = 2'b01;
		14'h1b54: color = 2'b01;
		14'h1b55: color = 2'b00;
		14'h1b56: color = 2'b01;
		14'h1b57: color = 2'b01;
		14'h1b58: color = 2'b01;
		14'h1b59: color = 2'b01;
		14'h1b5a: color = 2'b01;
		14'h1b5b: color = 2'b01;
		14'h1b5c: color = 2'b01;
		14'h1b5d: color = 2'b01;
		14'h1b5e: color = 2'b01;
		14'h1b5f: color = 2'b00;
		14'h1b60: color = 2'b00;
		14'h1b61: color = 2'b01;
		14'h1b62: color = 2'b00;
		14'h1b63: color = 2'b01;
		14'h1b64: color = 2'b11;
		14'h1b65: color = 2'b11;
		14'h1b66: color = 2'b11;
		14'h1b67: color = 2'b11;
		14'h1b68: color = 2'b11;
		14'h1b69: color = 2'b11;
		14'h1b6a: color = 2'b11;
		14'h1b6b: color = 2'b11;
		14'h1b6c: color = 2'b11;
		14'h1b6d: color = 2'b11;
		14'h1b6e: color = 2'b11;
		14'h1b6f: color = 2'b11;
		14'h1b70: color = 2'b11;
		14'h1b71: color = 2'b11;
		14'h1b72: color = 2'b11;
		14'h1b73: color = 2'b11;
		14'h1b74: color = 2'b11;
		14'h1b75: color = 2'b11;
		14'h1b76: color = 2'b11;
		14'h1b77: color = 2'b11;
		14'h1b78: color = 2'b11;
		14'h1b79: color = 2'b11;
		14'h1b7a: color = 2'b11;
		14'h1b7b: color = 2'b11;
		14'h1b7c: color = 2'b11;
		14'h1b7d: color = 2'b11;
		14'h1b7e: color = 2'b11;
		14'h1b7f: color = 2'b11;
		14'h1b80: color = 2'b11;
		14'h1b81: color = 2'b11;
		14'h1b82: color = 2'b11;
		14'h1b83: color = 2'b11;
		14'h1b84: color = 2'b11;
		14'h1b85: color = 2'b11;
		14'h1b86: color = 2'b11;
		14'h1b87: color = 2'b11;
		14'h1b88: color = 2'b11;
		14'h1b89: color = 2'b11;
		14'h1b8a: color = 2'b11;
		14'h1b8b: color = 2'b11;
		14'h1b8c: color = 2'b11;
		14'h1b8d: color = 2'b11;
		14'h1b8e: color = 2'b11;
		14'h1b8f: color = 2'b11;
		14'h1b90: color = 2'b11;
		14'h1b91: color = 2'b11;
		14'h1b92: color = 2'b11;
		14'h1b93: color = 2'b11;
		14'h1b94: color = 2'b11;
		14'h1b95: color = 2'b11;
		14'h1b96: color = 2'b11;
		14'h1b97: color = 2'b11;
		14'h1b98: color = 2'b11;
		14'h1b99: color = 2'b11;
		14'h1b9a: color = 2'b11;
		14'h1b9b: color = 2'b11;
		14'h1b9c: color = 2'b11;
		14'h1b9d: color = 2'b11;
		14'h1b9e: color = 2'b11;
		14'h1b9f: color = 2'b11;
		14'h1ba0: color = 2'b11;
		14'h1ba1: color = 2'b11;
		14'h1ba2: color = 2'b10;
		14'h1ba3: color = 2'b10;
		14'h1ba4: color = 2'b10;
		14'h1ba5: color = 2'b11;
		14'h1ba6: color = 2'b10;
		14'h1ba7: color = 2'b10;
		14'h1ba8: color = 2'b10;
		14'h1ba9: color = 2'b01;
		14'h1baa: color = 2'b01;
		14'h1bab: color = 2'b01;
		14'h1bac: color = 2'b00;
		14'h1bad: color = 2'b01;
		14'h1bae: color = 2'b01;
		14'h1baf: color = 2'b01;
		14'h1bb0: color = 2'b11;
		14'h1bb1: color = 2'b11;
		14'h1bb2: color = 2'b11;
		14'h1bb3: color = 2'b11;
		14'h1bb4: color = 2'b11;
		14'h1bb5: color = 2'b11;
		14'h1bb6: color = 2'b11;
		14'h1bb7: color = 2'b10;
		14'h1bb8: color = 2'b10;
		14'h1bb9: color = 2'b11;
		14'h1bba: color = 2'b10;
		14'h1bbb: color = 2'b10;
		14'h1bbc: color = 2'b10;
		14'h1bbd: color = 2'b11;
		14'h1bbe: color = 2'b10;
		14'h1bbf: color = 2'b10;
		14'h1bc0: color = 2'b10;
		14'h1bc1: color = 2'b10;
		14'h1bc2: color = 2'b10;
		14'h1bc3: color = 2'b10;
		14'h1bc4: color = 2'b01;
		14'h1bc5: color = 2'b01;
		14'h1bc6: color = 2'b01;
		14'h1bc7: color = 2'b01;
		14'h1bc8: color = 2'b01;
		14'h1bc9: color = 2'b10;
		14'h1bca: color = 2'b01;
		14'h1bcb: color = 2'b01;
		14'h1bcc: color = 2'b10;
		14'h1bcd: color = 2'b11;
		14'h1bce: color = 2'b11;
		14'h1bcf: color = 2'b10;
		14'h1bd0: color = 2'b01;
		14'h1bd1: color = 2'b00;
		14'h1bd2: color = 2'b01;
		14'h1bd3: color = 2'b01;
		14'h1bd4: color = 2'b01;
		14'h1bd5: color = 2'b01;
		14'h1bd6: color = 2'b01;
		14'h1bd7: color = 2'b01;
		14'h1bd8: color = 2'b01;
		14'h1bd9: color = 2'b01;
		14'h1bda: color = 2'b01;
		14'h1bdb: color = 2'b01;
		14'h1bdc: color = 2'b01;
		14'h1bdd: color = 2'b01;
		14'h1bde: color = 2'b01;
		14'h1bdf: color = 2'b01;
		14'h1be0: color = 2'b00;
		14'h1be1: color = 2'b00;
		14'h1be2: color = 2'b00;
		14'h1be3: color = 2'b10;
		14'h1be4: color = 2'b11;
		14'h1be5: color = 2'b11;
		14'h1be6: color = 2'b11;
		14'h1be7: color = 2'b11;
		14'h1be8: color = 2'b11;
		14'h1be9: color = 2'b11;
		14'h1bea: color = 2'b11;
		14'h1beb: color = 2'b11;
		14'h1bec: color = 2'b11;
		14'h1bed: color = 2'b11;
		14'h1bee: color = 2'b11;
		14'h1bef: color = 2'b11;
		14'h1bf0: color = 2'b11;
		14'h1bf1: color = 2'b11;
		14'h1bf2: color = 2'b11;
		14'h1bf3: color = 2'b11;
		14'h1bf4: color = 2'b11;
		14'h1bf5: color = 2'b11;
		14'h1bf6: color = 2'b11;
		14'h1bf7: color = 2'b11;
		14'h1bf8: color = 2'b11;
		14'h1bf9: color = 2'b11;
		14'h1bfa: color = 2'b11;
		14'h1bfb: color = 2'b11;
		14'h1bfc: color = 2'b11;
		14'h1bfd: color = 2'b11;
		14'h1bfe: color = 2'b11;
		14'h1bff: color = 2'b11;
		14'h1c00: color = 2'b11;
		14'h1c01: color = 2'b11;
		14'h1c02: color = 2'b11;
		14'h1c03: color = 2'b11;
		14'h1c04: color = 2'b11;
		14'h1c05: color = 2'b11;
		14'h1c06: color = 2'b11;
		14'h1c07: color = 2'b11;
		14'h1c08: color = 2'b11;
		14'h1c09: color = 2'b11;
		14'h1c0a: color = 2'b11;
		14'h1c0b: color = 2'b11;
		14'h1c0c: color = 2'b11;
		14'h1c0d: color = 2'b11;
		14'h1c0e: color = 2'b11;
		14'h1c0f: color = 2'b11;
		14'h1c10: color = 2'b11;
		14'h1c11: color = 2'b11;
		14'h1c12: color = 2'b11;
		14'h1c13: color = 2'b11;
		14'h1c14: color = 2'b11;
		14'h1c15: color = 2'b11;
		14'h1c16: color = 2'b11;
		14'h1c17: color = 2'b11;
		14'h1c18: color = 2'b11;
		14'h1c19: color = 2'b11;
		14'h1c1a: color = 2'b11;
		14'h1c1b: color = 2'b11;
		14'h1c1c: color = 2'b11;
		14'h1c1d: color = 2'b11;
		14'h1c1e: color = 2'b11;
		14'h1c1f: color = 2'b11;
		14'h1c20: color = 2'b11;
		14'h1c21: color = 2'b11;
		14'h1c22: color = 2'b10;
		14'h1c23: color = 2'b10;
		14'h1c24: color = 2'b10;
		14'h1c25: color = 2'b11;
		14'h1c26: color = 2'b10;
		14'h1c27: color = 2'b10;
		14'h1c28: color = 2'b10;
		14'h1c29: color = 2'b01;
		14'h1c2a: color = 2'b01;
		14'h1c2b: color = 2'b01;
		14'h1c2c: color = 2'b00;
		14'h1c2d: color = 2'b01;
		14'h1c2e: color = 2'b01;
		14'h1c2f: color = 2'b01;
		14'h1c30: color = 2'b11;
		14'h1c31: color = 2'b11;
		14'h1c32: color = 2'b11;
		14'h1c33: color = 2'b11;
		14'h1c34: color = 2'b11;
		14'h1c35: color = 2'b11;
		14'h1c36: color = 2'b11;
		14'h1c37: color = 2'b10;
		14'h1c38: color = 2'b10;
		14'h1c39: color = 2'b11;
		14'h1c3a: color = 2'b10;
		14'h1c3b: color = 2'b10;
		14'h1c3c: color = 2'b10;
		14'h1c3d: color = 2'b11;
		14'h1c3e: color = 2'b10;
		14'h1c3f: color = 2'b10;
		14'h1c40: color = 2'b10;
		14'h1c41: color = 2'b10;
		14'h1c42: color = 2'b10;
		14'h1c43: color = 2'b10;
		14'h1c44: color = 2'b01;
		14'h1c45: color = 2'b01;
		14'h1c46: color = 2'b01;
		14'h1c47: color = 2'b01;
		14'h1c48: color = 2'b01;
		14'h1c49: color = 2'b10;
		14'h1c4a: color = 2'b01;
		14'h1c4b: color = 2'b01;
		14'h1c4c: color = 2'b10;
		14'h1c4d: color = 2'b11;
		14'h1c4e: color = 2'b11;
		14'h1c4f: color = 2'b10;
		14'h1c50: color = 2'b01;
		14'h1c51: color = 2'b00;
		14'h1c52: color = 2'b01;
		14'h1c53: color = 2'b01;
		14'h1c54: color = 2'b01;
		14'h1c55: color = 2'b01;
		14'h1c56: color = 2'b01;
		14'h1c57: color = 2'b01;
		14'h1c58: color = 2'b01;
		14'h1c59: color = 2'b01;
		14'h1c5a: color = 2'b01;
		14'h1c5b: color = 2'b01;
		14'h1c5c: color = 2'b01;
		14'h1c5d: color = 2'b01;
		14'h1c5e: color = 2'b01;
		14'h1c5f: color = 2'b01;
		14'h1c60: color = 2'b00;
		14'h1c61: color = 2'b00;
		14'h1c62: color = 2'b00;
		14'h1c63: color = 2'b10;
		14'h1c64: color = 2'b11;
		14'h1c65: color = 2'b11;
		14'h1c66: color = 2'b11;
		14'h1c67: color = 2'b11;
		14'h1c68: color = 2'b11;
		14'h1c69: color = 2'b11;
		14'h1c6a: color = 2'b11;
		14'h1c6b: color = 2'b11;
		14'h1c6c: color = 2'b11;
		14'h1c6d: color = 2'b11;
		14'h1c6e: color = 2'b11;
		14'h1c6f: color = 2'b11;
		14'h1c70: color = 2'b11;
		14'h1c71: color = 2'b11;
		14'h1c72: color = 2'b11;
		14'h1c73: color = 2'b11;
		14'h1c74: color = 2'b11;
		14'h1c75: color = 2'b11;
		14'h1c76: color = 2'b11;
		14'h1c77: color = 2'b11;
		14'h1c78: color = 2'b11;
		14'h1c79: color = 2'b11;
		14'h1c7a: color = 2'b11;
		14'h1c7b: color = 2'b11;
		14'h1c7c: color = 2'b11;
		14'h1c7d: color = 2'b11;
		14'h1c7e: color = 2'b11;
		14'h1c7f: color = 2'b11;
		14'h1c80: color = 2'b11;
		14'h1c81: color = 2'b11;
		14'h1c82: color = 2'b11;
		14'h1c83: color = 2'b11;
		14'h1c84: color = 2'b11;
		14'h1c85: color = 2'b11;
		14'h1c86: color = 2'b11;
		14'h1c87: color = 2'b11;
		14'h1c88: color = 2'b11;
		14'h1c89: color = 2'b11;
		14'h1c8a: color = 2'b11;
		14'h1c8b: color = 2'b11;
		14'h1c8c: color = 2'b11;
		14'h1c8d: color = 2'b11;
		14'h1c8e: color = 2'b11;
		14'h1c8f: color = 2'b11;
		14'h1c90: color = 2'b11;
		14'h1c91: color = 2'b11;
		14'h1c92: color = 2'b11;
		14'h1c93: color = 2'b11;
		14'h1c94: color = 2'b11;
		14'h1c95: color = 2'b11;
		14'h1c96: color = 2'b11;
		14'h1c97: color = 2'b11;
		14'h1c98: color = 2'b11;
		14'h1c99: color = 2'b11;
		14'h1c9a: color = 2'b11;
		14'h1c9b: color = 2'b11;
		14'h1c9c: color = 2'b11;
		14'h1c9d: color = 2'b11;
		14'h1c9e: color = 2'b11;
		14'h1c9f: color = 2'b11;
		14'h1ca0: color = 2'b11;
		14'h1ca1: color = 2'b11;
		14'h1ca2: color = 2'b10;
		14'h1ca3: color = 2'b10;
		14'h1ca4: color = 2'b10;
		14'h1ca5: color = 2'b11;
		14'h1ca6: color = 2'b01;
		14'h1ca7: color = 2'b10;
		14'h1ca8: color = 2'b10;
		14'h1ca9: color = 2'b01;
		14'h1caa: color = 2'b01;
		14'h1cab: color = 2'b00;
		14'h1cac: color = 2'b00;
		14'h1cad: color = 2'b00;
		14'h1cae: color = 2'b01;
		14'h1caf: color = 2'b01;
		14'h1cb0: color = 2'b10;
		14'h1cb1: color = 2'b11;
		14'h1cb2: color = 2'b11;
		14'h1cb3: color = 2'b11;
		14'h1cb4: color = 2'b11;
		14'h1cb5: color = 2'b11;
		14'h1cb6: color = 2'b11;
		14'h1cb7: color = 2'b11;
		14'h1cb8: color = 2'b11;
		14'h1cb9: color = 2'b11;
		14'h1cba: color = 2'b10;
		14'h1cbb: color = 2'b11;
		14'h1cbc: color = 2'b10;
		14'h1cbd: color = 2'b10;
		14'h1cbe: color = 2'b10;
		14'h1cbf: color = 2'b10;
		14'h1cc0: color = 2'b10;
		14'h1cc1: color = 2'b10;
		14'h1cc2: color = 2'b01;
		14'h1cc3: color = 2'b01;
		14'h1cc4: color = 2'b01;
		14'h1cc5: color = 2'b01;
		14'h1cc6: color = 2'b10;
		14'h1cc7: color = 2'b10;
		14'h1cc8: color = 2'b10;
		14'h1cc9: color = 2'b10;
		14'h1cca: color = 2'b10;
		14'h1ccb: color = 2'b10;
		14'h1ccc: color = 2'b11;
		14'h1ccd: color = 2'b11;
		14'h1cce: color = 2'b10;
		14'h1ccf: color = 2'b10;
		14'h1cd0: color = 2'b01;
		14'h1cd1: color = 2'b01;
		14'h1cd2: color = 2'b01;
		14'h1cd3: color = 2'b01;
		14'h1cd4: color = 2'b01;
		14'h1cd5: color = 2'b01;
		14'h1cd6: color = 2'b01;
		14'h1cd7: color = 2'b01;
		14'h1cd8: color = 2'b01;
		14'h1cd9: color = 2'b01;
		14'h1cda: color = 2'b01;
		14'h1cdb: color = 2'b01;
		14'h1cdc: color = 2'b01;
		14'h1cdd: color = 2'b01;
		14'h1cde: color = 2'b10;
		14'h1cdf: color = 2'b01;
		14'h1ce0: color = 2'b00;
		14'h1ce1: color = 2'b00;
		14'h1ce2: color = 2'b00;
		14'h1ce3: color = 2'b01;
		14'h1ce4: color = 2'b11;
		14'h1ce5: color = 2'b11;
		14'h1ce6: color = 2'b11;
		14'h1ce7: color = 2'b11;
		14'h1ce8: color = 2'b11;
		14'h1ce9: color = 2'b11;
		14'h1cea: color = 2'b11;
		14'h1ceb: color = 2'b11;
		14'h1cec: color = 2'b11;
		14'h1ced: color = 2'b11;
		14'h1cee: color = 2'b11;
		14'h1cef: color = 2'b11;
		14'h1cf0: color = 2'b11;
		14'h1cf1: color = 2'b11;
		14'h1cf2: color = 2'b11;
		14'h1cf3: color = 2'b11;
		14'h1cf4: color = 2'b11;
		14'h1cf5: color = 2'b11;
		14'h1cf6: color = 2'b11;
		14'h1cf7: color = 2'b11;
		14'h1cf8: color = 2'b11;
		14'h1cf9: color = 2'b11;
		14'h1cfa: color = 2'b11;
		14'h1cfb: color = 2'b11;
		14'h1cfc: color = 2'b11;
		14'h1cfd: color = 2'b11;
		14'h1cfe: color = 2'b11;
		14'h1cff: color = 2'b11;
		14'h1d00: color = 2'b11;
		14'h1d01: color = 2'b11;
		14'h1d02: color = 2'b11;
		14'h1d03: color = 2'b11;
		14'h1d04: color = 2'b11;
		14'h1d05: color = 2'b11;
		14'h1d06: color = 2'b11;
		14'h1d07: color = 2'b11;
		14'h1d08: color = 2'b11;
		14'h1d09: color = 2'b11;
		14'h1d0a: color = 2'b11;
		14'h1d0b: color = 2'b11;
		14'h1d0c: color = 2'b11;
		14'h1d0d: color = 2'b11;
		14'h1d0e: color = 2'b11;
		14'h1d0f: color = 2'b11;
		14'h1d10: color = 2'b11;
		14'h1d11: color = 2'b11;
		14'h1d12: color = 2'b11;
		14'h1d13: color = 2'b11;
		14'h1d14: color = 2'b11;
		14'h1d15: color = 2'b11;
		14'h1d16: color = 2'b11;
		14'h1d17: color = 2'b11;
		14'h1d18: color = 2'b11;
		14'h1d19: color = 2'b11;
		14'h1d1a: color = 2'b11;
		14'h1d1b: color = 2'b11;
		14'h1d1c: color = 2'b11;
		14'h1d1d: color = 2'b11;
		14'h1d1e: color = 2'b11;
		14'h1d1f: color = 2'b11;
		14'h1d20: color = 2'b11;
		14'h1d21: color = 2'b11;
		14'h1d22: color = 2'b11;
		14'h1d23: color = 2'b10;
		14'h1d24: color = 2'b10;
		14'h1d25: color = 2'b11;
		14'h1d26: color = 2'b01;
		14'h1d27: color = 2'b00;
		14'h1d28: color = 2'b00;
		14'h1d29: color = 2'b01;
		14'h1d2a: color = 2'b01;
		14'h1d2b: color = 2'b00;
		14'h1d2c: color = 2'b01;
		14'h1d2d: color = 2'b01;
		14'h1d2e: color = 2'b01;
		14'h1d2f: color = 2'b10;
		14'h1d30: color = 2'b10;
		14'h1d31: color = 2'b11;
		14'h1d32: color = 2'b11;
		14'h1d33: color = 2'b11;
		14'h1d34: color = 2'b11;
		14'h1d35: color = 2'b11;
		14'h1d36: color = 2'b11;
		14'h1d37: color = 2'b11;
		14'h1d38: color = 2'b11;
		14'h1d39: color = 2'b11;
		14'h1d3a: color = 2'b11;
		14'h1d3b: color = 2'b11;
		14'h1d3c: color = 2'b10;
		14'h1d3d: color = 2'b10;
		14'h1d3e: color = 2'b10;
		14'h1d3f: color = 2'b10;
		14'h1d40: color = 2'b10;
		14'h1d41: color = 2'b10;
		14'h1d42: color = 2'b10;
		14'h1d43: color = 2'b10;
		14'h1d44: color = 2'b10;
		14'h1d45: color = 2'b10;
		14'h1d46: color = 2'b10;
		14'h1d47: color = 2'b10;
		14'h1d48: color = 2'b10;
		14'h1d49: color = 2'b10;
		14'h1d4a: color = 2'b10;
		14'h1d4b: color = 2'b10;
		14'h1d4c: color = 2'b11;
		14'h1d4d: color = 2'b11;
		14'h1d4e: color = 2'b11;
		14'h1d4f: color = 2'b10;
		14'h1d50: color = 2'b10;
		14'h1d51: color = 2'b01;
		14'h1d52: color = 2'b01;
		14'h1d53: color = 2'b10;
		14'h1d54: color = 2'b01;
		14'h1d55: color = 2'b01;
		14'h1d56: color = 2'b01;
		14'h1d57: color = 2'b01;
		14'h1d58: color = 2'b01;
		14'h1d59: color = 2'b01;
		14'h1d5a: color = 2'b01;
		14'h1d5b: color = 2'b01;
		14'h1d5c: color = 2'b10;
		14'h1d5d: color = 2'b10;
		14'h1d5e: color = 2'b01;
		14'h1d5f: color = 2'b01;
		14'h1d60: color = 2'b01;
		14'h1d61: color = 2'b00;
		14'h1d62: color = 2'b00;
		14'h1d63: color = 2'b10;
		14'h1d64: color = 2'b11;
		14'h1d65: color = 2'b11;
		14'h1d66: color = 2'b11;
		14'h1d67: color = 2'b11;
		14'h1d68: color = 2'b11;
		14'h1d69: color = 2'b11;
		14'h1d6a: color = 2'b11;
		14'h1d6b: color = 2'b11;
		14'h1d6c: color = 2'b11;
		14'h1d6d: color = 2'b11;
		14'h1d6e: color = 2'b11;
		14'h1d6f: color = 2'b11;
		14'h1d70: color = 2'b11;
		14'h1d71: color = 2'b11;
		14'h1d72: color = 2'b11;
		14'h1d73: color = 2'b11;
		14'h1d74: color = 2'b11;
		14'h1d75: color = 2'b11;
		14'h1d76: color = 2'b11;
		14'h1d77: color = 2'b11;
		14'h1d78: color = 2'b11;
		14'h1d79: color = 2'b11;
		14'h1d7a: color = 2'b11;
		14'h1d7b: color = 2'b11;
		14'h1d7c: color = 2'b11;
		14'h1d7d: color = 2'b11;
		14'h1d7e: color = 2'b11;
		14'h1d7f: color = 2'b11;
		14'h1d80: color = 2'b11;
		14'h1d81: color = 2'b11;
		14'h1d82: color = 2'b11;
		14'h1d83: color = 2'b11;
		14'h1d84: color = 2'b11;
		14'h1d85: color = 2'b11;
		14'h1d86: color = 2'b11;
		14'h1d87: color = 2'b11;
		14'h1d88: color = 2'b11;
		14'h1d89: color = 2'b11;
		14'h1d8a: color = 2'b11;
		14'h1d8b: color = 2'b11;
		14'h1d8c: color = 2'b11;
		14'h1d8d: color = 2'b11;
		14'h1d8e: color = 2'b11;
		14'h1d8f: color = 2'b11;
		14'h1d90: color = 2'b11;
		14'h1d91: color = 2'b11;
		14'h1d92: color = 2'b11;
		14'h1d93: color = 2'b11;
		14'h1d94: color = 2'b11;
		14'h1d95: color = 2'b11;
		14'h1d96: color = 2'b11;
		14'h1d97: color = 2'b11;
		14'h1d98: color = 2'b11;
		14'h1d99: color = 2'b11;
		14'h1d9a: color = 2'b11;
		14'h1d9b: color = 2'b11;
		14'h1d9c: color = 2'b11;
		14'h1d9d: color = 2'b11;
		14'h1d9e: color = 2'b11;
		14'h1d9f: color = 2'b11;
		14'h1da0: color = 2'b11;
		14'h1da1: color = 2'b11;
		14'h1da2: color = 2'b11;
		14'h1da3: color = 2'b10;
		14'h1da4: color = 2'b10;
		14'h1da5: color = 2'b11;
		14'h1da6: color = 2'b10;
		14'h1da7: color = 2'b01;
		14'h1da8: color = 2'b01;
		14'h1da9: color = 2'b01;
		14'h1daa: color = 2'b00;
		14'h1dab: color = 2'b01;
		14'h1dac: color = 2'b01;
		14'h1dad: color = 2'b01;
		14'h1dae: color = 2'b01;
		14'h1daf: color = 2'b01;
		14'h1db0: color = 2'b10;
		14'h1db1: color = 2'b11;
		14'h1db2: color = 2'b11;
		14'h1db3: color = 2'b11;
		14'h1db4: color = 2'b11;
		14'h1db5: color = 2'b11;
		14'h1db6: color = 2'b11;
		14'h1db7: color = 2'b11;
		14'h1db8: color = 2'b11;
		14'h1db9: color = 2'b11;
		14'h1dba: color = 2'b10;
		14'h1dbb: color = 2'b11;
		14'h1dbc: color = 2'b10;
		14'h1dbd: color = 2'b11;
		14'h1dbe: color = 2'b10;
		14'h1dbf: color = 2'b10;
		14'h1dc0: color = 2'b10;
		14'h1dc1: color = 2'b10;
		14'h1dc2: color = 2'b10;
		14'h1dc3: color = 2'b10;
		14'h1dc4: color = 2'b10;
		14'h1dc5: color = 2'b10;
		14'h1dc6: color = 2'b10;
		14'h1dc7: color = 2'b10;
		14'h1dc8: color = 2'b10;
		14'h1dc9: color = 2'b10;
		14'h1dca: color = 2'b10;
		14'h1dcb: color = 2'b11;
		14'h1dcc: color = 2'b11;
		14'h1dcd: color = 2'b11;
		14'h1dce: color = 2'b10;
		14'h1dcf: color = 2'b10;
		14'h1dd0: color = 2'b01;
		14'h1dd1: color = 2'b01;
		14'h1dd2: color = 2'b10;
		14'h1dd3: color = 2'b10;
		14'h1dd4: color = 2'b10;
		14'h1dd5: color = 2'b01;
		14'h1dd6: color = 2'b01;
		14'h1dd7: color = 2'b01;
		14'h1dd8: color = 2'b01;
		14'h1dd9: color = 2'b10;
		14'h1dda: color = 2'b01;
		14'h1ddb: color = 2'b10;
		14'h1ddc: color = 2'b01;
		14'h1ddd: color = 2'b10;
		14'h1dde: color = 2'b10;
		14'h1ddf: color = 2'b01;
		14'h1de0: color = 2'b01;
		14'h1de1: color = 2'b00;
		14'h1de2: color = 2'b00;
		14'h1de3: color = 2'b11;
		14'h1de4: color = 2'b11;
		14'h1de5: color = 2'b11;
		14'h1de6: color = 2'b11;
		14'h1de7: color = 2'b11;
		14'h1de8: color = 2'b11;
		14'h1de9: color = 2'b11;
		14'h1dea: color = 2'b11;
		14'h1deb: color = 2'b11;
		14'h1dec: color = 2'b11;
		14'h1ded: color = 2'b11;
		14'h1dee: color = 2'b11;
		14'h1def: color = 2'b11;
		14'h1df0: color = 2'b11;
		14'h1df1: color = 2'b11;
		14'h1df2: color = 2'b11;
		14'h1df3: color = 2'b11;
		14'h1df4: color = 2'b11;
		14'h1df5: color = 2'b11;
		14'h1df6: color = 2'b11;
		14'h1df7: color = 2'b11;
		14'h1df8: color = 2'b11;
		14'h1df9: color = 2'b11;
		14'h1dfa: color = 2'b11;
		14'h1dfb: color = 2'b11;
		14'h1dfc: color = 2'b11;
		14'h1dfd: color = 2'b11;
		14'h1dfe: color = 2'b11;
		14'h1dff: color = 2'b11;
		14'h1e00: color = 2'b11;
		14'h1e01: color = 2'b11;
		14'h1e02: color = 2'b11;
		14'h1e03: color = 2'b11;
		14'h1e04: color = 2'b11;
		14'h1e05: color = 2'b11;
		14'h1e06: color = 2'b11;
		14'h1e07: color = 2'b11;
		14'h1e08: color = 2'b11;
		14'h1e09: color = 2'b11;
		14'h1e0a: color = 2'b11;
		14'h1e0b: color = 2'b11;
		14'h1e0c: color = 2'b11;
		14'h1e0d: color = 2'b11;
		14'h1e0e: color = 2'b11;
		14'h1e0f: color = 2'b11;
		14'h1e10: color = 2'b11;
		14'h1e11: color = 2'b11;
		14'h1e12: color = 2'b11;
		14'h1e13: color = 2'b11;
		14'h1e14: color = 2'b11;
		14'h1e15: color = 2'b11;
		14'h1e16: color = 2'b11;
		14'h1e17: color = 2'b11;
		14'h1e18: color = 2'b11;
		14'h1e19: color = 2'b11;
		14'h1e1a: color = 2'b11;
		14'h1e1b: color = 2'b11;
		14'h1e1c: color = 2'b11;
		14'h1e1d: color = 2'b11;
		14'h1e1e: color = 2'b11;
		14'h1e1f: color = 2'b11;
		14'h1e20: color = 2'b11;
		14'h1e21: color = 2'b11;
		14'h1e22: color = 2'b11;
		14'h1e23: color = 2'b11;
		14'h1e24: color = 2'b00;
		14'h1e25: color = 2'b10;
		14'h1e26: color = 2'b11;
		14'h1e27: color = 2'b10;
		14'h1e28: color = 2'b10;
		14'h1e29: color = 2'b01;
		14'h1e2a: color = 2'b01;
		14'h1e2b: color = 2'b01;
		14'h1e2c: color = 2'b01;
		14'h1e2d: color = 2'b01;
		14'h1e2e: color = 2'b01;
		14'h1e2f: color = 2'b10;
		14'h1e30: color = 2'b10;
		14'h1e31: color = 2'b11;
		14'h1e32: color = 2'b11;
		14'h1e33: color = 2'b11;
		14'h1e34: color = 2'b11;
		14'h1e35: color = 2'b11;
		14'h1e36: color = 2'b11;
		14'h1e37: color = 2'b11;
		14'h1e38: color = 2'b11;
		14'h1e39: color = 2'b11;
		14'h1e3a: color = 2'b11;
		14'h1e3b: color = 2'b11;
		14'h1e3c: color = 2'b11;
		14'h1e3d: color = 2'b11;
		14'h1e3e: color = 2'b10;
		14'h1e3f: color = 2'b11;
		14'h1e40: color = 2'b10;
		14'h1e41: color = 2'b10;
		14'h1e42: color = 2'b10;
		14'h1e43: color = 2'b10;
		14'h1e44: color = 2'b10;
		14'h1e45: color = 2'b10;
		14'h1e46: color = 2'b10;
		14'h1e47: color = 2'b10;
		14'h1e48: color = 2'b10;
		14'h1e49: color = 2'b10;
		14'h1e4a: color = 2'b11;
		14'h1e4b: color = 2'b11;
		14'h1e4c: color = 2'b11;
		14'h1e4d: color = 2'b11;
		14'h1e4e: color = 2'b10;
		14'h1e4f: color = 2'b10;
		14'h1e50: color = 2'b01;
		14'h1e51: color = 2'b10;
		14'h1e52: color = 2'b01;
		14'h1e53: color = 2'b01;
		14'h1e54: color = 2'b10;
		14'h1e55: color = 2'b10;
		14'h1e56: color = 2'b10;
		14'h1e57: color = 2'b10;
		14'h1e58: color = 2'b10;
		14'h1e59: color = 2'b10;
		14'h1e5a: color = 2'b01;
		14'h1e5b: color = 2'b10;
		14'h1e5c: color = 2'b10;
		14'h1e5d: color = 2'b01;
		14'h1e5e: color = 2'b10;
		14'h1e5f: color = 2'b10;
		14'h1e60: color = 2'b00;
		14'h1e61: color = 2'b00;
		14'h1e62: color = 2'b00;
		14'h1e63: color = 2'b11;
		14'h1e64: color = 2'b11;
		14'h1e65: color = 2'b11;
		14'h1e66: color = 2'b11;
		14'h1e67: color = 2'b11;
		14'h1e68: color = 2'b11;
		14'h1e69: color = 2'b11;
		14'h1e6a: color = 2'b11;
		14'h1e6b: color = 2'b11;
		14'h1e6c: color = 2'b11;
		14'h1e6d: color = 2'b11;
		14'h1e6e: color = 2'b11;
		14'h1e6f: color = 2'b11;
		14'h1e70: color = 2'b11;
		14'h1e71: color = 2'b11;
		14'h1e72: color = 2'b11;
		14'h1e73: color = 2'b11;
		14'h1e74: color = 2'b11;
		14'h1e75: color = 2'b11;
		14'h1e76: color = 2'b11;
		14'h1e77: color = 2'b11;
		14'h1e78: color = 2'b11;
		14'h1e79: color = 2'b11;
		14'h1e7a: color = 2'b11;
		14'h1e7b: color = 2'b11;
		14'h1e7c: color = 2'b11;
		14'h1e7d: color = 2'b11;
		14'h1e7e: color = 2'b11;
		14'h1e7f: color = 2'b11;
		14'h1e80: color = 2'b11;
		14'h1e81: color = 2'b11;
		14'h1e82: color = 2'b11;
		14'h1e83: color = 2'b11;
		14'h1e84: color = 2'b11;
		14'h1e85: color = 2'b11;
		14'h1e86: color = 2'b11;
		14'h1e87: color = 2'b11;
		14'h1e88: color = 2'b11;
		14'h1e89: color = 2'b11;
		14'h1e8a: color = 2'b11;
		14'h1e8b: color = 2'b11;
		14'h1e8c: color = 2'b11;
		14'h1e8d: color = 2'b11;
		14'h1e8e: color = 2'b11;
		14'h1e8f: color = 2'b11;
		14'h1e90: color = 2'b11;
		14'h1e91: color = 2'b11;
		14'h1e92: color = 2'b11;
		14'h1e93: color = 2'b11;
		14'h1e94: color = 2'b11;
		14'h1e95: color = 2'b11;
		14'h1e96: color = 2'b11;
		14'h1e97: color = 2'b11;
		14'h1e98: color = 2'b11;
		14'h1e99: color = 2'b11;
		14'h1e9a: color = 2'b11;
		14'h1e9b: color = 2'b11;
		14'h1e9c: color = 2'b11;
		14'h1e9d: color = 2'b11;
		14'h1e9e: color = 2'b11;
		14'h1e9f: color = 2'b11;
		14'h1ea0: color = 2'b11;
		14'h1ea1: color = 2'b11;
		14'h1ea2: color = 2'b11;
		14'h1ea3: color = 2'b11;
		14'h1ea4: color = 2'b00;
		14'h1ea5: color = 2'b01;
		14'h1ea6: color = 2'b11;
		14'h1ea7: color = 2'b10;
		14'h1ea8: color = 2'b10;
		14'h1ea9: color = 2'b10;
		14'h1eaa: color = 2'b11;
		14'h1eab: color = 2'b10;
		14'h1eac: color = 2'b01;
		14'h1ead: color = 2'b01;
		14'h1eae: color = 2'b01;
		14'h1eaf: color = 2'b01;
		14'h1eb0: color = 2'b10;
		14'h1eb1: color = 2'b11;
		14'h1eb2: color = 2'b11;
		14'h1eb3: color = 2'b11;
		14'h1eb4: color = 2'b11;
		14'h1eb5: color = 2'b11;
		14'h1eb6: color = 2'b11;
		14'h1eb7: color = 2'b10;
		14'h1eb8: color = 2'b10;
		14'h1eb9: color = 2'b11;
		14'h1eba: color = 2'b10;
		14'h1ebb: color = 2'b10;
		14'h1ebc: color = 2'b10;
		14'h1ebd: color = 2'b10;
		14'h1ebe: color = 2'b10;
		14'h1ebf: color = 2'b10;
		14'h1ec0: color = 2'b10;
		14'h1ec1: color = 2'b10;
		14'h1ec2: color = 2'b10;
		14'h1ec3: color = 2'b10;
		14'h1ec4: color = 2'b10;
		14'h1ec5: color = 2'b10;
		14'h1ec6: color = 2'b10;
		14'h1ec7: color = 2'b11;
		14'h1ec8: color = 2'b11;
		14'h1ec9: color = 2'b11;
		14'h1eca: color = 2'b11;
		14'h1ecb: color = 2'b11;
		14'h1ecc: color = 2'b10;
		14'h1ecd: color = 2'b11;
		14'h1ece: color = 2'b10;
		14'h1ecf: color = 2'b10;
		14'h1ed0: color = 2'b10;
		14'h1ed1: color = 2'b01;
		14'h1ed2: color = 2'b10;
		14'h1ed3: color = 2'b10;
		14'h1ed4: color = 2'b10;
		14'h1ed5: color = 2'b10;
		14'h1ed6: color = 2'b10;
		14'h1ed7: color = 2'b10;
		14'h1ed8: color = 2'b10;
		14'h1ed9: color = 2'b01;
		14'h1eda: color = 2'b10;
		14'h1edb: color = 2'b10;
		14'h1edc: color = 2'b01;
		14'h1edd: color = 2'b10;
		14'h1ede: color = 2'b01;
		14'h1edf: color = 2'b01;
		14'h1ee0: color = 2'b00;
		14'h1ee1: color = 2'b00;
		14'h1ee2: color = 2'b10;
		14'h1ee3: color = 2'b11;
		14'h1ee4: color = 2'b11;
		14'h1ee5: color = 2'b11;
		14'h1ee6: color = 2'b11;
		14'h1ee7: color = 2'b11;
		14'h1ee8: color = 2'b11;
		14'h1ee9: color = 2'b11;
		14'h1eea: color = 2'b11;
		14'h1eeb: color = 2'b11;
		14'h1eec: color = 2'b11;
		14'h1eed: color = 2'b11;
		14'h1eee: color = 2'b11;
		14'h1eef: color = 2'b11;
		14'h1ef0: color = 2'b11;
		14'h1ef1: color = 2'b11;
		14'h1ef2: color = 2'b11;
		14'h1ef3: color = 2'b11;
		14'h1ef4: color = 2'b11;
		14'h1ef5: color = 2'b11;
		14'h1ef6: color = 2'b11;
		14'h1ef7: color = 2'b11;
		14'h1ef8: color = 2'b11;
		14'h1ef9: color = 2'b11;
		14'h1efa: color = 2'b11;
		14'h1efb: color = 2'b11;
		14'h1efc: color = 2'b11;
		14'h1efd: color = 2'b11;
		14'h1efe: color = 2'b11;
		14'h1eff: color = 2'b11;
		14'h1f00: color = 2'b11;
		14'h1f01: color = 2'b11;
		14'h1f02: color = 2'b11;
		14'h1f03: color = 2'b11;
		14'h1f04: color = 2'b11;
		14'h1f05: color = 2'b11;
		14'h1f06: color = 2'b11;
		14'h1f07: color = 2'b11;
		14'h1f08: color = 2'b11;
		14'h1f09: color = 2'b11;
		14'h1f0a: color = 2'b11;
		14'h1f0b: color = 2'b11;
		14'h1f0c: color = 2'b11;
		14'h1f0d: color = 2'b11;
		14'h1f0e: color = 2'b11;
		14'h1f0f: color = 2'b11;
		14'h1f10: color = 2'b11;
		14'h1f11: color = 2'b11;
		14'h1f12: color = 2'b11;
		14'h1f13: color = 2'b11;
		14'h1f14: color = 2'b11;
		14'h1f15: color = 2'b11;
		14'h1f16: color = 2'b11;
		14'h1f17: color = 2'b11;
		14'h1f18: color = 2'b11;
		14'h1f19: color = 2'b11;
		14'h1f1a: color = 2'b11;
		14'h1f1b: color = 2'b11;
		14'h1f1c: color = 2'b11;
		14'h1f1d: color = 2'b11;
		14'h1f1e: color = 2'b11;
		14'h1f1f: color = 2'b11;
		14'h1f20: color = 2'b11;
		14'h1f21: color = 2'b11;
		14'h1f22: color = 2'b11;
		14'h1f23: color = 2'b11;
		14'h1f24: color = 2'b11;
		14'h1f25: color = 2'b00;
		14'h1f26: color = 2'b01;
		14'h1f27: color = 2'b11;
		14'h1f28: color = 2'b11;
		14'h1f29: color = 2'b11;
		14'h1f2a: color = 2'b11;
		14'h1f2b: color = 2'b10;
		14'h1f2c: color = 2'b01;
		14'h1f2d: color = 2'b01;
		14'h1f2e: color = 2'b01;
		14'h1f2f: color = 2'b10;
		14'h1f30: color = 2'b10;
		14'h1f31: color = 2'b10;
		14'h1f32: color = 2'b11;
		14'h1f33: color = 2'b11;
		14'h1f34: color = 2'b10;
		14'h1f35: color = 2'b11;
		14'h1f36: color = 2'b11;
		14'h1f37: color = 2'b11;
		14'h1f38: color = 2'b11;
		14'h1f39: color = 2'b11;
		14'h1f3a: color = 2'b11;
		14'h1f3b: color = 2'b11;
		14'h1f3c: color = 2'b11;
		14'h1f3d: color = 2'b11;
		14'h1f3e: color = 2'b11;
		14'h1f3f: color = 2'b10;
		14'h1f40: color = 2'b11;
		14'h1f41: color = 2'b10;
		14'h1f42: color = 2'b10;
		14'h1f43: color = 2'b10;
		14'h1f44: color = 2'b10;
		14'h1f45: color = 2'b10;
		14'h1f46: color = 2'b10;
		14'h1f47: color = 2'b10;
		14'h1f48: color = 2'b10;
		14'h1f49: color = 2'b10;
		14'h1f4a: color = 2'b11;
		14'h1f4b: color = 2'b11;
		14'h1f4c: color = 2'b11;
		14'h1f4d: color = 2'b11;
		14'h1f4e: color = 2'b10;
		14'h1f4f: color = 2'b10;
		14'h1f50: color = 2'b01;
		14'h1f51: color = 2'b10;
		14'h1f52: color = 2'b01;
		14'h1f53: color = 2'b01;
		14'h1f54: color = 2'b10;
		14'h1f55: color = 2'b10;
		14'h1f56: color = 2'b01;
		14'h1f57: color = 2'b10;
		14'h1f58: color = 2'b10;
		14'h1f59: color = 2'b10;
		14'h1f5a: color = 2'b10;
		14'h1f5b: color = 2'b01;
		14'h1f5c: color = 2'b10;
		14'h1f5d: color = 2'b01;
		14'h1f5e: color = 2'b10;
		14'h1f5f: color = 2'b01;
		14'h1f60: color = 2'b00;
		14'h1f61: color = 2'b00;
		14'h1f62: color = 2'b11;
		14'h1f63: color = 2'b11;
		14'h1f64: color = 2'b11;
		14'h1f65: color = 2'b11;
		14'h1f66: color = 2'b11;
		14'h1f67: color = 2'b11;
		14'h1f68: color = 2'b11;
		14'h1f69: color = 2'b11;
		14'h1f6a: color = 2'b11;
		14'h1f6b: color = 2'b11;
		14'h1f6c: color = 2'b11;
		14'h1f6d: color = 2'b11;
		14'h1f6e: color = 2'b11;
		14'h1f6f: color = 2'b11;
		14'h1f70: color = 2'b11;
		14'h1f71: color = 2'b11;
		14'h1f72: color = 2'b11;
		14'h1f73: color = 2'b11;
		14'h1f74: color = 2'b11;
		14'h1f75: color = 2'b11;
		14'h1f76: color = 2'b11;
		14'h1f77: color = 2'b11;
		14'h1f78: color = 2'b11;
		14'h1f79: color = 2'b11;
		14'h1f7a: color = 2'b11;
		14'h1f7b: color = 2'b11;
		14'h1f7c: color = 2'b11;
		14'h1f7d: color = 2'b11;
		14'h1f7e: color = 2'b11;
		14'h1f7f: color = 2'b11;
		14'h1f80: color = 2'b11;
		14'h1f81: color = 2'b11;
		14'h1f82: color = 2'b11;
		14'h1f83: color = 2'b11;
		14'h1f84: color = 2'b11;
		14'h1f85: color = 2'b11;
		14'h1f86: color = 2'b11;
		14'h1f87: color = 2'b11;
		14'h1f88: color = 2'b11;
		14'h1f89: color = 2'b11;
		14'h1f8a: color = 2'b11;
		14'h1f8b: color = 2'b11;
		14'h1f8c: color = 2'b11;
		14'h1f8d: color = 2'b11;
		14'h1f8e: color = 2'b11;
		14'h1f8f: color = 2'b11;
		14'h1f90: color = 2'b11;
		14'h1f91: color = 2'b11;
		14'h1f92: color = 2'b11;
		14'h1f93: color = 2'b11;
		14'h1f94: color = 2'b11;
		14'h1f95: color = 2'b11;
		14'h1f96: color = 2'b11;
		14'h1f97: color = 2'b11;
		14'h1f98: color = 2'b11;
		14'h1f99: color = 2'b11;
		14'h1f9a: color = 2'b11;
		14'h1f9b: color = 2'b11;
		14'h1f9c: color = 2'b11;
		14'h1f9d: color = 2'b11;
		14'h1f9e: color = 2'b11;
		14'h1f9f: color = 2'b11;
		14'h1fa0: color = 2'b11;
		14'h1fa1: color = 2'b11;
		14'h1fa2: color = 2'b11;
		14'h1fa3: color = 2'b11;
		14'h1fa4: color = 2'b11;
		14'h1fa5: color = 2'b00;
		14'h1fa6: color = 2'b00;
		14'h1fa7: color = 2'b10;
		14'h1fa8: color = 2'b10;
		14'h1fa9: color = 2'b11;
		14'h1faa: color = 2'b11;
		14'h1fab: color = 2'b11;
		14'h1fac: color = 2'b10;
		14'h1fad: color = 2'b01;
		14'h1fae: color = 2'b01;
		14'h1faf: color = 2'b01;
		14'h1fb0: color = 2'b10;
		14'h1fb1: color = 2'b10;
		14'h1fb2: color = 2'b11;
		14'h1fb3: color = 2'b11;
		14'h1fb4: color = 2'b11;
		14'h1fb5: color = 2'b11;
		14'h1fb6: color = 2'b11;
		14'h1fb7: color = 2'b11;
		14'h1fb8: color = 2'b11;
		14'h1fb9: color = 2'b11;
		14'h1fba: color = 2'b11;
		14'h1fbb: color = 2'b11;
		14'h1fbc: color = 2'b11;
		14'h1fbd: color = 2'b10;
		14'h1fbe: color = 2'b11;
		14'h1fbf: color = 2'b10;
		14'h1fc0: color = 2'b11;
		14'h1fc1: color = 2'b10;
		14'h1fc2: color = 2'b11;
		14'h1fc3: color = 2'b10;
		14'h1fc4: color = 2'b10;
		14'h1fc5: color = 2'b10;
		14'h1fc6: color = 2'b10;
		14'h1fc7: color = 2'b11;
		14'h1fc8: color = 2'b11;
		14'h1fc9: color = 2'b10;
		14'h1fca: color = 2'b11;
		14'h1fcb: color = 2'b10;
		14'h1fcc: color = 2'b11;
		14'h1fcd: color = 2'b10;
		14'h1fce: color = 2'b10;
		14'h1fcf: color = 2'b10;
		14'h1fd0: color = 2'b10;
		14'h1fd1: color = 2'b01;
		14'h1fd2: color = 2'b01;
		14'h1fd3: color = 2'b10;
		14'h1fd4: color = 2'b10;
		14'h1fd5: color = 2'b10;
		14'h1fd6: color = 2'b10;
		14'h1fd7: color = 2'b10;
		14'h1fd8: color = 2'b10;
		14'h1fd9: color = 2'b10;
		14'h1fda: color = 2'b10;
		14'h1fdb: color = 2'b10;
		14'h1fdc: color = 2'b01;
		14'h1fdd: color = 2'b10;
		14'h1fde: color = 2'b01;
		14'h1fdf: color = 2'b01;
		14'h1fe0: color = 2'b00;
		14'h1fe1: color = 2'b00;
		14'h1fe2: color = 2'b11;
		14'h1fe3: color = 2'b11;
		14'h1fe4: color = 2'b11;
		14'h1fe5: color = 2'b11;
		14'h1fe6: color = 2'b11;
		14'h1fe7: color = 2'b11;
		14'h1fe8: color = 2'b11;
		14'h1fe9: color = 2'b11;
		14'h1fea: color = 2'b11;
		14'h1feb: color = 2'b11;
		14'h1fec: color = 2'b11;
		14'h1fed: color = 2'b11;
		14'h1fee: color = 2'b11;
		14'h1fef: color = 2'b11;
		14'h1ff0: color = 2'b11;
		14'h1ff1: color = 2'b11;
		14'h1ff2: color = 2'b11;
		14'h1ff3: color = 2'b11;
		14'h1ff4: color = 2'b11;
		14'h1ff5: color = 2'b11;
		14'h1ff6: color = 2'b11;
		14'h1ff7: color = 2'b11;
		14'h1ff8: color = 2'b11;
		14'h1ff9: color = 2'b11;
		14'h1ffa: color = 2'b11;
		14'h1ffb: color = 2'b11;
		14'h1ffc: color = 2'b11;
		14'h1ffd: color = 2'b11;
		14'h1ffe: color = 2'b11;
		14'h1fff: color = 2'b11;
		14'h2000: color = 2'b11;
		14'h2001: color = 2'b11;
		14'h2002: color = 2'b11;
		14'h2003: color = 2'b11;
		14'h2004: color = 2'b11;
		14'h2005: color = 2'b11;
		14'h2006: color = 2'b11;
		14'h2007: color = 2'b11;
		14'h2008: color = 2'b11;
		14'h2009: color = 2'b11;
		14'h200a: color = 2'b11;
		14'h200b: color = 2'b11;
		14'h200c: color = 2'b11;
		14'h200d: color = 2'b11;
		14'h200e: color = 2'b11;
		14'h200f: color = 2'b11;
		14'h2010: color = 2'b11;
		14'h2011: color = 2'b11;
		14'h2012: color = 2'b11;
		14'h2013: color = 2'b11;
		14'h2014: color = 2'b11;
		14'h2015: color = 2'b11;
		14'h2016: color = 2'b11;
		14'h2017: color = 2'b11;
		14'h2018: color = 2'b11;
		14'h2019: color = 2'b11;
		14'h201a: color = 2'b11;
		14'h201b: color = 2'b11;
		14'h201c: color = 2'b11;
		14'h201d: color = 2'b11;
		14'h201e: color = 2'b11;
		14'h201f: color = 2'b11;
		14'h2020: color = 2'b11;
		14'h2021: color = 2'b11;
		14'h2022: color = 2'b11;
		14'h2023: color = 2'b11;
		14'h2024: color = 2'b11;
		14'h2025: color = 2'b11;
		14'h2026: color = 2'b00;
		14'h2027: color = 2'b01;
		14'h2028: color = 2'b01;
		14'h2029: color = 2'b11;
		14'h202a: color = 2'b11;
		14'h202b: color = 2'b11;
		14'h202c: color = 2'b10;
		14'h202d: color = 2'b01;
		14'h202e: color = 2'b01;
		14'h202f: color = 2'b01;
		14'h2030: color = 2'b10;
		14'h2031: color = 2'b10;
		14'h2032: color = 2'b11;
		14'h2033: color = 2'b11;
		14'h2034: color = 2'b11;
		14'h2035: color = 2'b11;
		14'h2036: color = 2'b11;
		14'h2037: color = 2'b10;
		14'h2038: color = 2'b10;
		14'h2039: color = 2'b11;
		14'h203a: color = 2'b11;
		14'h203b: color = 2'b11;
		14'h203c: color = 2'b11;
		14'h203d: color = 2'b11;
		14'h203e: color = 2'b11;
		14'h203f: color = 2'b10;
		14'h2040: color = 2'b11;
		14'h2041: color = 2'b10;
		14'h2042: color = 2'b10;
		14'h2043: color = 2'b10;
		14'h2044: color = 2'b01;
		14'h2045: color = 2'b10;
		14'h2046: color = 2'b10;
		14'h2047: color = 2'b11;
		14'h2048: color = 2'b11;
		14'h2049: color = 2'b11;
		14'h204a: color = 2'b10;
		14'h204b: color = 2'b11;
		14'h204c: color = 2'b10;
		14'h204d: color = 2'b11;
		14'h204e: color = 2'b10;
		14'h204f: color = 2'b10;
		14'h2050: color = 2'b01;
		14'h2051: color = 2'b10;
		14'h2052: color = 2'b01;
		14'h2053: color = 2'b01;
		14'h2054: color = 2'b10;
		14'h2055: color = 2'b10;
		14'h2056: color = 2'b10;
		14'h2057: color = 2'b10;
		14'h2058: color = 2'b10;
		14'h2059: color = 2'b10;
		14'h205a: color = 2'b10;
		14'h205b: color = 2'b10;
		14'h205c: color = 2'b10;
		14'h205d: color = 2'b01;
		14'h205e: color = 2'b10;
		14'h205f: color = 2'b00;
		14'h2060: color = 2'b00;
		14'h2061: color = 2'b11;
		14'h2062: color = 2'b11;
		14'h2063: color = 2'b11;
		14'h2064: color = 2'b11;
		14'h2065: color = 2'b11;
		14'h2066: color = 2'b11;
		14'h2067: color = 2'b11;
		14'h2068: color = 2'b11;
		14'h2069: color = 2'b11;
		14'h206a: color = 2'b11;
		14'h206b: color = 2'b11;
		14'h206c: color = 2'b11;
		14'h206d: color = 2'b11;
		14'h206e: color = 2'b11;
		14'h206f: color = 2'b11;
		14'h2070: color = 2'b11;
		14'h2071: color = 2'b11;
		14'h2072: color = 2'b11;
		14'h2073: color = 2'b11;
		14'h2074: color = 2'b11;
		14'h2075: color = 2'b11;
		14'h2076: color = 2'b11;
		14'h2077: color = 2'b11;
		14'h2078: color = 2'b11;
		14'h2079: color = 2'b11;
		14'h207a: color = 2'b11;
		14'h207b: color = 2'b11;
		14'h207c: color = 2'b11;
		14'h207d: color = 2'b11;
		14'h207e: color = 2'b11;
		14'h207f: color = 2'b11;
		14'h2080: color = 2'b11;
		14'h2081: color = 2'b11;
		14'h2082: color = 2'b11;
		14'h2083: color = 2'b11;
		14'h2084: color = 2'b11;
		14'h2085: color = 2'b11;
		14'h2086: color = 2'b11;
		14'h2087: color = 2'b11;
		14'h2088: color = 2'b11;
		14'h2089: color = 2'b11;
		14'h208a: color = 2'b11;
		14'h208b: color = 2'b11;
		14'h208c: color = 2'b11;
		14'h208d: color = 2'b11;
		14'h208e: color = 2'b11;
		14'h208f: color = 2'b11;
		14'h2090: color = 2'b11;
		14'h2091: color = 2'b11;
		14'h2092: color = 2'b11;
		14'h2093: color = 2'b11;
		14'h2094: color = 2'b11;
		14'h2095: color = 2'b11;
		14'h2096: color = 2'b11;
		14'h2097: color = 2'b11;
		14'h2098: color = 2'b11;
		14'h2099: color = 2'b11;
		14'h209a: color = 2'b11;
		14'h209b: color = 2'b11;
		14'h209c: color = 2'b11;
		14'h209d: color = 2'b11;
		14'h209e: color = 2'b11;
		14'h209f: color = 2'b11;
		14'h20a0: color = 2'b11;
		14'h20a1: color = 2'b11;
		14'h20a2: color = 2'b11;
		14'h20a3: color = 2'b11;
		14'h20a4: color = 2'b11;
		14'h20a5: color = 2'b11;
		14'h20a6: color = 2'b00;
		14'h20a7: color = 2'b00;
		14'h20a8: color = 2'b00;
		14'h20a9: color = 2'b10;
		14'h20aa: color = 2'b11;
		14'h20ab: color = 2'b11;
		14'h20ac: color = 2'b10;
		14'h20ad: color = 2'b01;
		14'h20ae: color = 2'b01;
		14'h20af: color = 2'b01;
		14'h20b0: color = 2'b10;
		14'h20b1: color = 2'b01;
		14'h20b2: color = 2'b11;
		14'h20b3: color = 2'b11;
		14'h20b4: color = 2'b11;
		14'h20b5: color = 2'b10;
		14'h20b6: color = 2'b11;
		14'h20b7: color = 2'b11;
		14'h20b8: color = 2'b11;
		14'h20b9: color = 2'b11;
		14'h20ba: color = 2'b10;
		14'h20bb: color = 2'b11;
		14'h20bc: color = 2'b11;
		14'h20bd: color = 2'b10;
		14'h20be: color = 2'b11;
		14'h20bf: color = 2'b10;
		14'h20c0: color = 2'b10;
		14'h20c1: color = 2'b10;
		14'h20c2: color = 2'b10;
		14'h20c3: color = 2'b10;
		14'h20c4: color = 2'b01;
		14'h20c5: color = 2'b10;
		14'h20c6: color = 2'b11;
		14'h20c7: color = 2'b11;
		14'h20c8: color = 2'b11;
		14'h20c9: color = 2'b10;
		14'h20ca: color = 2'b11;
		14'h20cb: color = 2'b11;
		14'h20cc: color = 2'b11;
		14'h20cd: color = 2'b11;
		14'h20ce: color = 2'b10;
		14'h20cf: color = 2'b10;
		14'h20d0: color = 2'b10;
		14'h20d1: color = 2'b10;
		14'h20d2: color = 2'b01;
		14'h20d3: color = 2'b01;
		14'h20d4: color = 2'b01;
		14'h20d5: color = 2'b10;
		14'h20d6: color = 2'b10;
		14'h20d7: color = 2'b10;
		14'h20d8: color = 2'b10;
		14'h20d9: color = 2'b10;
		14'h20da: color = 2'b10;
		14'h20db: color = 2'b10;
		14'h20dc: color = 2'b01;
		14'h20dd: color = 2'b01;
		14'h20de: color = 2'b01;
		14'h20df: color = 2'b00;
		14'h20e0: color = 2'b00;
		14'h20e1: color = 2'b11;
		14'h20e2: color = 2'b11;
		14'h20e3: color = 2'b11;
		14'h20e4: color = 2'b11;
		14'h20e5: color = 2'b11;
		14'h20e6: color = 2'b11;
		14'h20e7: color = 2'b11;
		14'h20e8: color = 2'b11;
		14'h20e9: color = 2'b11;
		14'h20ea: color = 2'b11;
		14'h20eb: color = 2'b11;
		14'h20ec: color = 2'b11;
		14'h20ed: color = 2'b11;
		14'h20ee: color = 2'b11;
		14'h20ef: color = 2'b11;
		14'h20f0: color = 2'b11;
		14'h20f1: color = 2'b11;
		14'h20f2: color = 2'b11;
		14'h20f3: color = 2'b11;
		14'h20f4: color = 2'b11;
		14'h20f5: color = 2'b11;
		14'h20f6: color = 2'b11;
		14'h20f7: color = 2'b11;
		14'h20f8: color = 2'b11;
		14'h20f9: color = 2'b11;
		14'h20fa: color = 2'b11;
		14'h20fb: color = 2'b11;
		14'h20fc: color = 2'b11;
		14'h20fd: color = 2'b11;
		14'h20fe: color = 2'b11;
		14'h20ff: color = 2'b11;
		14'h2100: color = 2'b11;
		14'h2101: color = 2'b11;
		14'h2102: color = 2'b11;
		14'h2103: color = 2'b11;
		14'h2104: color = 2'b11;
		14'h2105: color = 2'b11;
		14'h2106: color = 2'b11;
		14'h2107: color = 2'b11;
		14'h2108: color = 2'b11;
		14'h2109: color = 2'b11;
		14'h210a: color = 2'b11;
		14'h210b: color = 2'b11;
		14'h210c: color = 2'b11;
		14'h210d: color = 2'b11;
		14'h210e: color = 2'b11;
		14'h210f: color = 2'b11;
		14'h2110: color = 2'b11;
		14'h2111: color = 2'b11;
		14'h2112: color = 2'b11;
		14'h2113: color = 2'b11;
		14'h2114: color = 2'b11;
		14'h2115: color = 2'b11;
		14'h2116: color = 2'b11;
		14'h2117: color = 2'b11;
		14'h2118: color = 2'b11;
		14'h2119: color = 2'b11;
		14'h211a: color = 2'b11;
		14'h211b: color = 2'b11;
		14'h211c: color = 2'b11;
		14'h211d: color = 2'b11;
		14'h211e: color = 2'b11;
		14'h211f: color = 2'b11;
		14'h2120: color = 2'b11;
		14'h2121: color = 2'b11;
		14'h2122: color = 2'b11;
		14'h2123: color = 2'b11;
		14'h2124: color = 2'b11;
		14'h2125: color = 2'b10;
		14'h2126: color = 2'b00;
		14'h2127: color = 2'b00;
		14'h2128: color = 2'b00;
		14'h2129: color = 2'b10;
		14'h212a: color = 2'b10;
		14'h212b: color = 2'b11;
		14'h212c: color = 2'b10;
		14'h212d: color = 2'b10;
		14'h212e: color = 2'b01;
		14'h212f: color = 2'b10;
		14'h2130: color = 2'b01;
		14'h2131: color = 2'b10;
		14'h2132: color = 2'b10;
		14'h2133: color = 2'b11;
		14'h2134: color = 2'b11;
		14'h2135: color = 2'b11;
		14'h2136: color = 2'b11;
		14'h2137: color = 2'b10;
		14'h2138: color = 2'b10;
		14'h2139: color = 2'b11;
		14'h213a: color = 2'b11;
		14'h213b: color = 2'b11;
		14'h213c: color = 2'b10;
		14'h213d: color = 2'b11;
		14'h213e: color = 2'b10;
		14'h213f: color = 2'b11;
		14'h2140: color = 2'b10;
		14'h2141: color = 2'b10;
		14'h2142: color = 2'b10;
		14'h2143: color = 2'b01;
		14'h2144: color = 2'b01;
		14'h2145: color = 2'b01;
		14'h2146: color = 2'b11;
		14'h2147: color = 2'b11;
		14'h2148: color = 2'b11;
		14'h2149: color = 2'b11;
		14'h214a: color = 2'b11;
		14'h214b: color = 2'b11;
		14'h214c: color = 2'b11;
		14'h214d: color = 2'b11;
		14'h214e: color = 2'b11;
		14'h214f: color = 2'b10;
		14'h2150: color = 2'b10;
		14'h2151: color = 2'b01;
		14'h2152: color = 2'b10;
		14'h2153: color = 2'b01;
		14'h2154: color = 2'b01;
		14'h2155: color = 2'b01;
		14'h2156: color = 2'b01;
		14'h2157: color = 2'b10;
		14'h2158: color = 2'b10;
		14'h2159: color = 2'b10;
		14'h215a: color = 2'b01;
		14'h215b: color = 2'b10;
		14'h215c: color = 2'b10;
		14'h215d: color = 2'b01;
		14'h215e: color = 2'b01;
		14'h215f: color = 2'b00;
		14'h2160: color = 2'b01;
		14'h2161: color = 2'b11;
		14'h2162: color = 2'b11;
		14'h2163: color = 2'b11;
		14'h2164: color = 2'b11;
		14'h2165: color = 2'b11;
		14'h2166: color = 2'b11;
		14'h2167: color = 2'b11;
		14'h2168: color = 2'b11;
		14'h2169: color = 2'b11;
		14'h216a: color = 2'b11;
		14'h216b: color = 2'b11;
		14'h216c: color = 2'b11;
		14'h216d: color = 2'b11;
		14'h216e: color = 2'b11;
		14'h216f: color = 2'b11;
		14'h2170: color = 2'b11;
		14'h2171: color = 2'b11;
		14'h2172: color = 2'b11;
		14'h2173: color = 2'b11;
		14'h2174: color = 2'b11;
		14'h2175: color = 2'b11;
		14'h2176: color = 2'b11;
		14'h2177: color = 2'b11;
		14'h2178: color = 2'b11;
		14'h2179: color = 2'b11;
		14'h217a: color = 2'b11;
		14'h217b: color = 2'b11;
		14'h217c: color = 2'b11;
		14'h217d: color = 2'b11;
		14'h217e: color = 2'b11;
		14'h217f: color = 2'b11;
		14'h2180: color = 2'b11;
		14'h2181: color = 2'b11;
		14'h2182: color = 2'b11;
		14'h2183: color = 2'b11;
		14'h2184: color = 2'b11;
		14'h2185: color = 2'b11;
		14'h2186: color = 2'b11;
		14'h2187: color = 2'b11;
		14'h2188: color = 2'b11;
		14'h2189: color = 2'b11;
		14'h218a: color = 2'b11;
		14'h218b: color = 2'b11;
		14'h218c: color = 2'b11;
		14'h218d: color = 2'b11;
		14'h218e: color = 2'b11;
		14'h218f: color = 2'b11;
		14'h2190: color = 2'b11;
		14'h2191: color = 2'b11;
		14'h2192: color = 2'b11;
		14'h2193: color = 2'b11;
		14'h2194: color = 2'b11;
		14'h2195: color = 2'b11;
		14'h2196: color = 2'b11;
		14'h2197: color = 2'b11;
		14'h2198: color = 2'b11;
		14'h2199: color = 2'b11;
		14'h219a: color = 2'b11;
		14'h219b: color = 2'b11;
		14'h219c: color = 2'b11;
		14'h219d: color = 2'b11;
		14'h219e: color = 2'b11;
		14'h219f: color = 2'b11;
		14'h21a0: color = 2'b11;
		14'h21a1: color = 2'b11;
		14'h21a2: color = 2'b11;
		14'h21a3: color = 2'b11;
		14'h21a4: color = 2'b11;
		14'h21a5: color = 2'b01;
		14'h21a6: color = 2'b01;
		14'h21a7: color = 2'b00;
		14'h21a8: color = 2'b00;
		14'h21a9: color = 2'b01;
		14'h21aa: color = 2'b10;
		14'h21ab: color = 2'b11;
		14'h21ac: color = 2'b10;
		14'h21ad: color = 2'b01;
		14'h21ae: color = 2'b01;
		14'h21af: color = 2'b10;
		14'h21b0: color = 2'b10;
		14'h21b1: color = 2'b10;
		14'h21b2: color = 2'b10;
		14'h21b3: color = 2'b11;
		14'h21b4: color = 2'b11;
		14'h21b5: color = 2'b10;
		14'h21b6: color = 2'b11;
		14'h21b7: color = 2'b11;
		14'h21b8: color = 2'b11;
		14'h21b9: color = 2'b11;
		14'h21ba: color = 2'b10;
		14'h21bb: color = 2'b11;
		14'h21bc: color = 2'b11;
		14'h21bd: color = 2'b10;
		14'h21be: color = 2'b10;
		14'h21bf: color = 2'b10;
		14'h21c0: color = 2'b10;
		14'h21c1: color = 2'b10;
		14'h21c2: color = 2'b01;
		14'h21c3: color = 2'b01;
		14'h21c4: color = 2'b01;
		14'h21c5: color = 2'b10;
		14'h21c6: color = 2'b10;
		14'h21c7: color = 2'b10;
		14'h21c8: color = 2'b10;
		14'h21c9: color = 2'b10;
		14'h21ca: color = 2'b10;
		14'h21cb: color = 2'b10;
		14'h21cc: color = 2'b11;
		14'h21cd: color = 2'b11;
		14'h21ce: color = 2'b10;
		14'h21cf: color = 2'b10;
		14'h21d0: color = 2'b01;
		14'h21d1: color = 2'b01;
		14'h21d2: color = 2'b01;
		14'h21d3: color = 2'b01;
		14'h21d4: color = 2'b01;
		14'h21d5: color = 2'b01;
		14'h21d6: color = 2'b01;
		14'h21d7: color = 2'b10;
		14'h21d8: color = 2'b10;
		14'h21d9: color = 2'b01;
		14'h21da: color = 2'b10;
		14'h21db: color = 2'b01;
		14'h21dc: color = 2'b01;
		14'h21dd: color = 2'b01;
		14'h21de: color = 2'b01;
		14'h21df: color = 2'b00;
		14'h21e0: color = 2'b11;
		14'h21e1: color = 2'b11;
		14'h21e2: color = 2'b11;
		14'h21e3: color = 2'b11;
		14'h21e4: color = 2'b11;
		14'h21e5: color = 2'b11;
		14'h21e6: color = 2'b11;
		14'h21e7: color = 2'b11;
		14'h21e8: color = 2'b11;
		14'h21e9: color = 2'b11;
		14'h21ea: color = 2'b11;
		14'h21eb: color = 2'b11;
		14'h21ec: color = 2'b11;
		14'h21ed: color = 2'b11;
		14'h21ee: color = 2'b11;
		14'h21ef: color = 2'b11;
		14'h21f0: color = 2'b11;
		14'h21f1: color = 2'b11;
		14'h21f2: color = 2'b11;
		14'h21f3: color = 2'b11;
		14'h21f4: color = 2'b11;
		14'h21f5: color = 2'b11;
		14'h21f6: color = 2'b11;
		14'h21f7: color = 2'b11;
		14'h21f8: color = 2'b11;
		14'h21f9: color = 2'b11;
		14'h21fa: color = 2'b11;
		14'h21fb: color = 2'b11;
		14'h21fc: color = 2'b11;
		14'h21fd: color = 2'b11;
		14'h21fe: color = 2'b11;
		14'h21ff: color = 2'b11;
		14'h2200: color = 2'b11;
		14'h2201: color = 2'b11;
		14'h2202: color = 2'b11;
		14'h2203: color = 2'b11;
		14'h2204: color = 2'b11;
		14'h2205: color = 2'b11;
		14'h2206: color = 2'b11;
		14'h2207: color = 2'b11;
		14'h2208: color = 2'b11;
		14'h2209: color = 2'b11;
		14'h220a: color = 2'b11;
		14'h220b: color = 2'b11;
		14'h220c: color = 2'b11;
		14'h220d: color = 2'b11;
		14'h220e: color = 2'b11;
		14'h220f: color = 2'b11;
		14'h2210: color = 2'b11;
		14'h2211: color = 2'b11;
		14'h2212: color = 2'b11;
		14'h2213: color = 2'b11;
		14'h2214: color = 2'b11;
		14'h2215: color = 2'b11;
		14'h2216: color = 2'b11;
		14'h2217: color = 2'b11;
		14'h2218: color = 2'b11;
		14'h2219: color = 2'b11;
		14'h221a: color = 2'b11;
		14'h221b: color = 2'b11;
		14'h221c: color = 2'b11;
		14'h221d: color = 2'b11;
		14'h221e: color = 2'b11;
		14'h221f: color = 2'b11;
		14'h2220: color = 2'b11;
		14'h2221: color = 2'b11;
		14'h2222: color = 2'b11;
		14'h2223: color = 2'b11;
		14'h2224: color = 2'b11;
		14'h2225: color = 2'b11;
		14'h2226: color = 2'b00;
		14'h2227: color = 2'b00;
		14'h2228: color = 2'b00;
		14'h2229: color = 2'b10;
		14'h222a: color = 2'b10;
		14'h222b: color = 2'b10;
		14'h222c: color = 2'b10;
		14'h222d: color = 2'b01;
		14'h222e: color = 2'b01;
		14'h222f: color = 2'b10;
		14'h2230: color = 2'b01;
		14'h2231: color = 2'b10;
		14'h2232: color = 2'b10;
		14'h2233: color = 2'b10;
		14'h2234: color = 2'b11;
		14'h2235: color = 2'b11;
		14'h2236: color = 2'b11;
		14'h2237: color = 2'b10;
		14'h2238: color = 2'b10;
		14'h2239: color = 2'b11;
		14'h223a: color = 2'b11;
		14'h223b: color = 2'b11;
		14'h223c: color = 2'b11;
		14'h223d: color = 2'b11;
		14'h223e: color = 2'b10;
		14'h223f: color = 2'b10;
		14'h2240: color = 2'b10;
		14'h2241: color = 2'b01;
		14'h2242: color = 2'b01;
		14'h2243: color = 2'b10;
		14'h2244: color = 2'b10;
		14'h2245: color = 2'b10;
		14'h2246: color = 2'b01;
		14'h2247: color = 2'b01;
		14'h2248: color = 2'b01;
		14'h2249: color = 2'b00;
		14'h224a: color = 2'b01;
		14'h224b: color = 2'b01;
		14'h224c: color = 2'b10;
		14'h224d: color = 2'b10;
		14'h224e: color = 2'b01;
		14'h224f: color = 2'b01;
		14'h2250: color = 2'b01;
		14'h2251: color = 2'b00;
		14'h2252: color = 2'b00;
		14'h2253: color = 2'b01;
		14'h2254: color = 2'b01;
		14'h2255: color = 2'b00;
		14'h2256: color = 2'b01;
		14'h2257: color = 2'b01;
		14'h2258: color = 2'b01;
		14'h2259: color = 2'b01;
		14'h225a: color = 2'b01;
		14'h225b: color = 2'b10;
		14'h225c: color = 2'b01;
		14'h225d: color = 2'b01;
		14'h225e: color = 2'b00;
		14'h225f: color = 2'b00;
		14'h2260: color = 2'b11;
		14'h2261: color = 2'b11;
		14'h2262: color = 2'b11;
		14'h2263: color = 2'b11;
		14'h2264: color = 2'b11;
		14'h2265: color = 2'b11;
		14'h2266: color = 2'b11;
		14'h2267: color = 2'b11;
		14'h2268: color = 2'b11;
		14'h2269: color = 2'b11;
		14'h226a: color = 2'b11;
		14'h226b: color = 2'b11;
		14'h226c: color = 2'b11;
		14'h226d: color = 2'b11;
		14'h226e: color = 2'b11;
		14'h226f: color = 2'b11;
		14'h2270: color = 2'b11;
		14'h2271: color = 2'b11;
		14'h2272: color = 2'b11;
		14'h2273: color = 2'b11;
		14'h2274: color = 2'b11;
		14'h2275: color = 2'b11;
		14'h2276: color = 2'b11;
		14'h2277: color = 2'b11;
		14'h2278: color = 2'b11;
		14'h2279: color = 2'b11;
		14'h227a: color = 2'b11;
		14'h227b: color = 2'b11;
		14'h227c: color = 2'b11;
		14'h227d: color = 2'b11;
		14'h227e: color = 2'b11;
		14'h227f: color = 2'b11;
		14'h2280: color = 2'b11;
		14'h2281: color = 2'b11;
		14'h2282: color = 2'b11;
		14'h2283: color = 2'b11;
		14'h2284: color = 2'b11;
		14'h2285: color = 2'b11;
		14'h2286: color = 2'b11;
		14'h2287: color = 2'b11;
		14'h2288: color = 2'b11;
		14'h2289: color = 2'b11;
		14'h228a: color = 2'b11;
		14'h228b: color = 2'b11;
		14'h228c: color = 2'b11;
		14'h228d: color = 2'b11;
		14'h228e: color = 2'b11;
		14'h228f: color = 2'b11;
		14'h2290: color = 2'b11;
		14'h2291: color = 2'b11;
		14'h2292: color = 2'b11;
		14'h2293: color = 2'b11;
		14'h2294: color = 2'b11;
		14'h2295: color = 2'b11;
		14'h2296: color = 2'b11;
		14'h2297: color = 2'b11;
		14'h2298: color = 2'b11;
		14'h2299: color = 2'b11;
		14'h229a: color = 2'b11;
		14'h229b: color = 2'b11;
		14'h229c: color = 2'b11;
		14'h229d: color = 2'b11;
		14'h229e: color = 2'b11;
		14'h229f: color = 2'b11;
		14'h22a0: color = 2'b11;
		14'h22a1: color = 2'b11;
		14'h22a2: color = 2'b11;
		14'h22a3: color = 2'b11;
		14'h22a4: color = 2'b11;
		14'h22a5: color = 2'b11;
		14'h22a6: color = 2'b00;
		14'h22a7: color = 2'b00;
		14'h22a8: color = 2'b00;
		14'h22a9: color = 2'b01;
		14'h22aa: color = 2'b10;
		14'h22ab: color = 2'b11;
		14'h22ac: color = 2'b10;
		14'h22ad: color = 2'b01;
		14'h22ae: color = 2'b01;
		14'h22af: color = 2'b10;
		14'h22b0: color = 2'b01;
		14'h22b1: color = 2'b10;
		14'h22b2: color = 2'b01;
		14'h22b3: color = 2'b10;
		14'h22b4: color = 2'b10;
		14'h22b5: color = 2'b11;
		14'h22b6: color = 2'b11;
		14'h22b7: color = 2'b10;
		14'h22b8: color = 2'b10;
		14'h22b9: color = 2'b11;
		14'h22ba: color = 2'b10;
		14'h22bb: color = 2'b11;
		14'h22bc: color = 2'b10;
		14'h22bd: color = 2'b10;
		14'h22be: color = 2'b10;
		14'h22bf: color = 2'b10;
		14'h22c0: color = 2'b01;
		14'h22c1: color = 2'b01;
		14'h22c2: color = 2'b10;
		14'h22c3: color = 2'b01;
		14'h22c4: color = 2'b01;
		14'h22c5: color = 2'b01;
		14'h22c6: color = 2'b01;
		14'h22c7: color = 2'b00;
		14'h22c8: color = 2'b00;
		14'h22c9: color = 2'b00;
		14'h22ca: color = 2'b00;
		14'h22cb: color = 2'b00;
		14'h22cc: color = 2'b00;
		14'h22cd: color = 2'b01;
		14'h22ce: color = 2'b00;
		14'h22cf: color = 2'b00;
		14'h22d0: color = 2'b00;
		14'h22d1: color = 2'b00;
		14'h22d2: color = 2'b00;
		14'h22d3: color = 2'b00;
		14'h22d4: color = 2'b00;
		14'h22d5: color = 2'b00;
		14'h22d6: color = 2'b01;
		14'h22d7: color = 2'b01;
		14'h22d8: color = 2'b01;
		14'h22d9: color = 2'b01;
		14'h22da: color = 2'b01;
		14'h22db: color = 2'b01;
		14'h22dc: color = 2'b01;
		14'h22dd: color = 2'b01;
		14'h22de: color = 2'b00;
		14'h22df: color = 2'b00;
		14'h22e0: color = 2'b11;
		14'h22e1: color = 2'b11;
		14'h22e2: color = 2'b11;
		14'h22e3: color = 2'b11;
		14'h22e4: color = 2'b11;
		14'h22e5: color = 2'b11;
		14'h22e6: color = 2'b11;
		14'h22e7: color = 2'b11;
		14'h22e8: color = 2'b11;
		14'h22e9: color = 2'b11;
		14'h22ea: color = 2'b11;
		14'h22eb: color = 2'b11;
		14'h22ec: color = 2'b11;
		14'h22ed: color = 2'b11;
		14'h22ee: color = 2'b11;
		14'h22ef: color = 2'b11;
		14'h22f0: color = 2'b11;
		14'h22f1: color = 2'b11;
		14'h22f2: color = 2'b11;
		14'h22f3: color = 2'b11;
		14'h22f4: color = 2'b11;
		14'h22f5: color = 2'b11;
		14'h22f6: color = 2'b11;
		14'h22f7: color = 2'b11;
		14'h22f8: color = 2'b11;
		14'h22f9: color = 2'b11;
		14'h22fa: color = 2'b11;
		14'h22fb: color = 2'b11;
		14'h22fc: color = 2'b11;
		14'h22fd: color = 2'b11;
		14'h22fe: color = 2'b11;
		14'h22ff: color = 2'b11;
		14'h2300: color = 2'b11;
		14'h2301: color = 2'b11;
		14'h2302: color = 2'b11;
		14'h2303: color = 2'b11;
		14'h2304: color = 2'b11;
		14'h2305: color = 2'b11;
		14'h2306: color = 2'b11;
		14'h2307: color = 2'b11;
		14'h2308: color = 2'b11;
		14'h2309: color = 2'b11;
		14'h230a: color = 2'b11;
		14'h230b: color = 2'b11;
		14'h230c: color = 2'b11;
		14'h230d: color = 2'b11;
		14'h230e: color = 2'b11;
		14'h230f: color = 2'b11;
		14'h2310: color = 2'b11;
		14'h2311: color = 2'b11;
		14'h2312: color = 2'b11;
		14'h2313: color = 2'b11;
		14'h2314: color = 2'b11;
		14'h2315: color = 2'b11;
		14'h2316: color = 2'b11;
		14'h2317: color = 2'b11;
		14'h2318: color = 2'b11;
		14'h2319: color = 2'b11;
		14'h231a: color = 2'b11;
		14'h231b: color = 2'b11;
		14'h231c: color = 2'b11;
		14'h231d: color = 2'b11;
		14'h231e: color = 2'b11;
		14'h231f: color = 2'b11;
		14'h2320: color = 2'b11;
		14'h2321: color = 2'b11;
		14'h2322: color = 2'b11;
		14'h2323: color = 2'b11;
		14'h2324: color = 2'b11;
		14'h2325: color = 2'b11;
		14'h2326: color = 2'b10;
		14'h2327: color = 2'b01;
		14'h2328: color = 2'b01;
		14'h2329: color = 2'b01;
		14'h232a: color = 2'b11;
		14'h232b: color = 2'b10;
		14'h232c: color = 2'b11;
		14'h232d: color = 2'b01;
		14'h232e: color = 2'b01;
		14'h232f: color = 2'b10;
		14'h2330: color = 2'b01;
		14'h2331: color = 2'b10;
		14'h2332: color = 2'b01;
		14'h2333: color = 2'b10;
		14'h2334: color = 2'b10;
		14'h2335: color = 2'b10;
		14'h2336: color = 2'b11;
		14'h2337: color = 2'b10;
		14'h2338: color = 2'b10;
		14'h2339: color = 2'b11;
		14'h233a: color = 2'b11;
		14'h233b: color = 2'b11;
		14'h233c: color = 2'b11;
		14'h233d: color = 2'b10;
		14'h233e: color = 2'b10;
		14'h233f: color = 2'b01;
		14'h2340: color = 2'b01;
		14'h2341: color = 2'b01;
		14'h2342: color = 2'b01;
		14'h2343: color = 2'b01;
		14'h2344: color = 2'b01;
		14'h2345: color = 2'b00;
		14'h2346: color = 2'b00;
		14'h2347: color = 2'b00;
		14'h2348: color = 2'b00;
		14'h2349: color = 2'b00;
		14'h234a: color = 2'b00;
		14'h234b: color = 2'b00;
		14'h234c: color = 2'b00;
		14'h234d: color = 2'b00;
		14'h234e: color = 2'b00;
		14'h234f: color = 2'b00;
		14'h2350: color = 2'b00;
		14'h2351: color = 2'b00;
		14'h2352: color = 2'b00;
		14'h2353: color = 2'b00;
		14'h2354: color = 2'b00;
		14'h2355: color = 2'b00;
		14'h2356: color = 2'b00;
		14'h2357: color = 2'b00;
		14'h2358: color = 2'b00;
		14'h2359: color = 2'b01;
		14'h235a: color = 2'b01;
		14'h235b: color = 2'b01;
		14'h235c: color = 2'b01;
		14'h235d: color = 2'b01;
		14'h235e: color = 2'b00;
		14'h235f: color = 2'b01;
		14'h2360: color = 2'b11;
		14'h2361: color = 2'b11;
		14'h2362: color = 2'b11;
		14'h2363: color = 2'b11;
		14'h2364: color = 2'b11;
		14'h2365: color = 2'b11;
		14'h2366: color = 2'b11;
		14'h2367: color = 2'b11;
		14'h2368: color = 2'b11;
		14'h2369: color = 2'b11;
		14'h236a: color = 2'b11;
		14'h236b: color = 2'b11;
		14'h236c: color = 2'b11;
		14'h236d: color = 2'b11;
		14'h236e: color = 2'b11;
		14'h236f: color = 2'b11;
		14'h2370: color = 2'b11;
		14'h2371: color = 2'b11;
		14'h2372: color = 2'b11;
		14'h2373: color = 2'b11;
		14'h2374: color = 2'b11;
		14'h2375: color = 2'b11;
		14'h2376: color = 2'b11;
		14'h2377: color = 2'b11;
		14'h2378: color = 2'b11;
		14'h2379: color = 2'b11;
		14'h237a: color = 2'b11;
		14'h237b: color = 2'b11;
		14'h237c: color = 2'b11;
		14'h237d: color = 2'b11;
		14'h237e: color = 2'b11;
		14'h237f: color = 2'b11;
		14'h2380: color = 2'b11;
		14'h2381: color = 2'b11;
		14'h2382: color = 2'b11;
		14'h2383: color = 2'b11;
		14'h2384: color = 2'b11;
		14'h2385: color = 2'b11;
		14'h2386: color = 2'b11;
		14'h2387: color = 2'b11;
		14'h2388: color = 2'b11;
		14'h2389: color = 2'b11;
		14'h238a: color = 2'b11;
		14'h238b: color = 2'b11;
		14'h238c: color = 2'b11;
		14'h238d: color = 2'b11;
		14'h238e: color = 2'b11;
		14'h238f: color = 2'b11;
		14'h2390: color = 2'b11;
		14'h2391: color = 2'b11;
		14'h2392: color = 2'b11;
		14'h2393: color = 2'b11;
		14'h2394: color = 2'b11;
		14'h2395: color = 2'b11;
		14'h2396: color = 2'b11;
		14'h2397: color = 2'b11;
		14'h2398: color = 2'b11;
		14'h2399: color = 2'b11;
		14'h239a: color = 2'b11;
		14'h239b: color = 2'b11;
		14'h239c: color = 2'b11;
		14'h239d: color = 2'b11;
		14'h239e: color = 2'b11;
		14'h239f: color = 2'b11;
		14'h23a0: color = 2'b11;
		14'h23a1: color = 2'b11;
		14'h23a2: color = 2'b11;
		14'h23a3: color = 2'b11;
		14'h23a4: color = 2'b11;
		14'h23a5: color = 2'b11;
		14'h23a6: color = 2'b10;
		14'h23a7: color = 2'b01;
		14'h23a8: color = 2'b01;
		14'h23a9: color = 2'b01;
		14'h23aa: color = 2'b10;
		14'h23ab: color = 2'b10;
		14'h23ac: color = 2'b10;
		14'h23ad: color = 2'b10;
		14'h23ae: color = 2'b01;
		14'h23af: color = 2'b01;
		14'h23b0: color = 2'b10;
		14'h23b1: color = 2'b01;
		14'h23b2: color = 2'b01;
		14'h23b3: color = 2'b10;
		14'h23b4: color = 2'b01;
		14'h23b5: color = 2'b10;
		14'h23b6: color = 2'b10;
		14'h23b7: color = 2'b10;
		14'h23b8: color = 2'b10;
		14'h23b9: color = 2'b11;
		14'h23ba: color = 2'b11;
		14'h23bb: color = 2'b11;
		14'h23bc: color = 2'b10;
		14'h23bd: color = 2'b10;
		14'h23be: color = 2'b00;
		14'h23bf: color = 2'b01;
		14'h23c0: color = 2'b01;
		14'h23c1: color = 2'b00;
		14'h23c2: color = 2'b00;
		14'h23c3: color = 2'b01;
		14'h23c4: color = 2'b00;
		14'h23c5: color = 2'b00;
		14'h23c6: color = 2'b00;
		14'h23c7: color = 2'b00;
		14'h23c8: color = 2'b00;
		14'h23c9: color = 2'b00;
		14'h23ca: color = 2'b00;
		14'h23cb: color = 2'b00;
		14'h23cc: color = 2'b00;
		14'h23cd: color = 2'b00;
		14'h23ce: color = 2'b00;
		14'h23cf: color = 2'b00;
		14'h23d0: color = 2'b00;
		14'h23d1: color = 2'b00;
		14'h23d2: color = 2'b00;
		14'h23d3: color = 2'b00;
		14'h23d4: color = 2'b00;
		14'h23d5: color = 2'b00;
		14'h23d6: color = 2'b00;
		14'h23d7: color = 2'b00;
		14'h23d8: color = 2'b00;
		14'h23d9: color = 2'b01;
		14'h23da: color = 2'b01;
		14'h23db: color = 2'b01;
		14'h23dc: color = 2'b01;
		14'h23dd: color = 2'b00;
		14'h23de: color = 2'b00;
		14'h23df: color = 2'b11;
		14'h23e0: color = 2'b11;
		14'h23e1: color = 2'b11;
		14'h23e2: color = 2'b11;
		14'h23e3: color = 2'b11;
		14'h23e4: color = 2'b11;
		14'h23e5: color = 2'b11;
		14'h23e6: color = 2'b11;
		14'h23e7: color = 2'b11;
		14'h23e8: color = 2'b11;
		14'h23e9: color = 2'b11;
		14'h23ea: color = 2'b11;
		14'h23eb: color = 2'b11;
		14'h23ec: color = 2'b11;
		14'h23ed: color = 2'b11;
		14'h23ee: color = 2'b11;
		14'h23ef: color = 2'b11;
		14'h23f0: color = 2'b11;
		14'h23f1: color = 2'b11;
		14'h23f2: color = 2'b11;
		14'h23f3: color = 2'b11;
		14'h23f4: color = 2'b11;
		14'h23f5: color = 2'b11;
		14'h23f6: color = 2'b11;
		14'h23f7: color = 2'b11;
		14'h23f8: color = 2'b11;
		14'h23f9: color = 2'b11;
		14'h23fa: color = 2'b11;
		14'h23fb: color = 2'b11;
		14'h23fc: color = 2'b11;
		14'h23fd: color = 2'b11;
		14'h23fe: color = 2'b11;
		14'h23ff: color = 2'b11;
		14'h2400: color = 2'b11;
		14'h2401: color = 2'b11;
		14'h2402: color = 2'b11;
		14'h2403: color = 2'b11;
		14'h2404: color = 2'b11;
		14'h2405: color = 2'b11;
		14'h2406: color = 2'b11;
		14'h2407: color = 2'b11;
		14'h2408: color = 2'b11;
		14'h2409: color = 2'b11;
		14'h240a: color = 2'b11;
		14'h240b: color = 2'b11;
		14'h240c: color = 2'b11;
		14'h240d: color = 2'b11;
		14'h240e: color = 2'b11;
		14'h240f: color = 2'b11;
		14'h2410: color = 2'b11;
		14'h2411: color = 2'b11;
		14'h2412: color = 2'b11;
		14'h2413: color = 2'b11;
		14'h2414: color = 2'b11;
		14'h2415: color = 2'b11;
		14'h2416: color = 2'b11;
		14'h2417: color = 2'b11;
		14'h2418: color = 2'b11;
		14'h2419: color = 2'b11;
		14'h241a: color = 2'b11;
		14'h241b: color = 2'b11;
		14'h241c: color = 2'b11;
		14'h241d: color = 2'b11;
		14'h241e: color = 2'b11;
		14'h241f: color = 2'b11;
		14'h2420: color = 2'b11;
		14'h2421: color = 2'b11;
		14'h2422: color = 2'b11;
		14'h2423: color = 2'b11;
		14'h2424: color = 2'b11;
		14'h2425: color = 2'b11;
		14'h2426: color = 2'b10;
		14'h2427: color = 2'b01;
		14'h2428: color = 2'b01;
		14'h2429: color = 2'b01;
		14'h242a: color = 2'b10;
		14'h242b: color = 2'b10;
		14'h242c: color = 2'b10;
		14'h242d: color = 2'b10;
		14'h242e: color = 2'b01;
		14'h242f: color = 2'b01;
		14'h2430: color = 2'b10;
		14'h2431: color = 2'b01;
		14'h2432: color = 2'b01;
		14'h2433: color = 2'b10;
		14'h2434: color = 2'b01;
		14'h2435: color = 2'b10;
		14'h2436: color = 2'b10;
		14'h2437: color = 2'b10;
		14'h2438: color = 2'b10;
		14'h2439: color = 2'b11;
		14'h243a: color = 2'b11;
		14'h243b: color = 2'b11;
		14'h243c: color = 2'b10;
		14'h243d: color = 2'b10;
		14'h243e: color = 2'b00;
		14'h243f: color = 2'b01;
		14'h2440: color = 2'b01;
		14'h2441: color = 2'b00;
		14'h2442: color = 2'b00;
		14'h2443: color = 2'b01;
		14'h2444: color = 2'b00;
		14'h2445: color = 2'b00;
		14'h2446: color = 2'b00;
		14'h2447: color = 2'b00;
		14'h2448: color = 2'b00;
		14'h2449: color = 2'b00;
		14'h244a: color = 2'b00;
		14'h244b: color = 2'b00;
		14'h244c: color = 2'b00;
		14'h244d: color = 2'b00;
		14'h244e: color = 2'b00;
		14'h244f: color = 2'b00;
		14'h2450: color = 2'b00;
		14'h2451: color = 2'b00;
		14'h2452: color = 2'b00;
		14'h2453: color = 2'b00;
		14'h2454: color = 2'b00;
		14'h2455: color = 2'b00;
		14'h2456: color = 2'b00;
		14'h2457: color = 2'b00;
		14'h2458: color = 2'b00;
		14'h2459: color = 2'b01;
		14'h245a: color = 2'b01;
		14'h245b: color = 2'b01;
		14'h245c: color = 2'b01;
		14'h245d: color = 2'b00;
		14'h245e: color = 2'b00;
		14'h245f: color = 2'b11;
		14'h2460: color = 2'b11;
		14'h2461: color = 2'b11;
		14'h2462: color = 2'b11;
		14'h2463: color = 2'b11;
		14'h2464: color = 2'b11;
		14'h2465: color = 2'b11;
		14'h2466: color = 2'b11;
		14'h2467: color = 2'b11;
		14'h2468: color = 2'b11;
		14'h2469: color = 2'b11;
		14'h246a: color = 2'b11;
		14'h246b: color = 2'b11;
		14'h246c: color = 2'b11;
		14'h246d: color = 2'b11;
		14'h246e: color = 2'b11;
		14'h246f: color = 2'b11;
		14'h2470: color = 2'b11;
		14'h2471: color = 2'b11;
		14'h2472: color = 2'b11;
		14'h2473: color = 2'b11;
		14'h2474: color = 2'b11;
		14'h2475: color = 2'b11;
		14'h2476: color = 2'b11;
		14'h2477: color = 2'b11;
		14'h2478: color = 2'b11;
		14'h2479: color = 2'b11;
		14'h247a: color = 2'b11;
		14'h247b: color = 2'b11;
		14'h247c: color = 2'b11;
		14'h247d: color = 2'b11;
		14'h247e: color = 2'b11;
		14'h247f: color = 2'b11;
		14'h2480: color = 2'b11;
		14'h2481: color = 2'b11;
		14'h2482: color = 2'b11;
		14'h2483: color = 2'b11;
		14'h2484: color = 2'b11;
		14'h2485: color = 2'b11;
		14'h2486: color = 2'b11;
		14'h2487: color = 2'b11;
		14'h2488: color = 2'b11;
		14'h2489: color = 2'b11;
		14'h248a: color = 2'b11;
		14'h248b: color = 2'b11;
		14'h248c: color = 2'b11;
		14'h248d: color = 2'b11;
		14'h248e: color = 2'b11;
		14'h248f: color = 2'b11;
		14'h2490: color = 2'b11;
		14'h2491: color = 2'b11;
		14'h2492: color = 2'b11;
		14'h2493: color = 2'b11;
		14'h2494: color = 2'b11;
		14'h2495: color = 2'b11;
		14'h2496: color = 2'b11;
		14'h2497: color = 2'b11;
		14'h2498: color = 2'b11;
		14'h2499: color = 2'b11;
		14'h249a: color = 2'b11;
		14'h249b: color = 2'b11;
		14'h249c: color = 2'b11;
		14'h249d: color = 2'b11;
		14'h249e: color = 2'b11;
		14'h249f: color = 2'b11;
		14'h24a0: color = 2'b11;
		14'h24a1: color = 2'b11;
		14'h24a2: color = 2'b11;
		14'h24a3: color = 2'b11;
		14'h24a4: color = 2'b11;
		14'h24a5: color = 2'b11;
		14'h24a6: color = 2'b11;
		14'h24a7: color = 2'b00;
		14'h24a8: color = 2'b00;
		14'h24a9: color = 2'b01;
		14'h24aa: color = 2'b10;
		14'h24ab: color = 2'b11;
		14'h24ac: color = 2'b10;
		14'h24ad: color = 2'b10;
		14'h24ae: color = 2'b01;
		14'h24af: color = 2'b10;
		14'h24b0: color = 2'b10;
		14'h24b1: color = 2'b01;
		14'h24b2: color = 2'b01;
		14'h24b3: color = 2'b01;
		14'h24b4: color = 2'b01;
		14'h24b5: color = 2'b01;
		14'h24b6: color = 2'b10;
		14'h24b7: color = 2'b10;
		14'h24b8: color = 2'b10;
		14'h24b9: color = 2'b11;
		14'h24ba: color = 2'b11;
		14'h24bb: color = 2'b11;
		14'h24bc: color = 2'b10;
		14'h24bd: color = 2'b00;
		14'h24be: color = 2'b01;
		14'h24bf: color = 2'b00;
		14'h24c0: color = 2'b00;
		14'h24c1: color = 2'b00;
		14'h24c2: color = 2'b00;
		14'h24c3: color = 2'b00;
		14'h24c4: color = 2'b00;
		14'h24c5: color = 2'b00;
		14'h24c6: color = 2'b00;
		14'h24c7: color = 2'b00;
		14'h24c8: color = 2'b00;
		14'h24c9: color = 2'b00;
		14'h24ca: color = 2'b00;
		14'h24cb: color = 2'b00;
		14'h24cc: color = 2'b00;
		14'h24cd: color = 2'b00;
		14'h24ce: color = 2'b00;
		14'h24cf: color = 2'b00;
		14'h24d0: color = 2'b00;
		14'h24d1: color = 2'b00;
		14'h24d2: color = 2'b00;
		14'h24d3: color = 2'b00;
		14'h24d4: color = 2'b00;
		14'h24d5: color = 2'b00;
		14'h24d6: color = 2'b00;
		14'h24d7: color = 2'b00;
		14'h24d8: color = 2'b00;
		14'h24d9: color = 2'b01;
		14'h24da: color = 2'b01;
		14'h24db: color = 2'b01;
		14'h24dc: color = 2'b01;
		14'h24dd: color = 2'b00;
		14'h24de: color = 2'b00;
		14'h24df: color = 2'b11;
		14'h24e0: color = 2'b11;
		14'h24e1: color = 2'b11;
		14'h24e2: color = 2'b11;
		14'h24e3: color = 2'b11;
		14'h24e4: color = 2'b11;
		14'h24e5: color = 2'b11;
		14'h24e6: color = 2'b11;
		14'h24e7: color = 2'b11;
		14'h24e8: color = 2'b11;
		14'h24e9: color = 2'b11;
		14'h24ea: color = 2'b11;
		14'h24eb: color = 2'b11;
		14'h24ec: color = 2'b11;
		14'h24ed: color = 2'b11;
		14'h24ee: color = 2'b11;
		14'h24ef: color = 2'b11;
		14'h24f0: color = 2'b11;
		14'h24f1: color = 2'b11;
		14'h24f2: color = 2'b11;
		14'h24f3: color = 2'b11;
		14'h24f4: color = 2'b11;
		14'h24f5: color = 2'b11;
		14'h24f6: color = 2'b11;
		14'h24f7: color = 2'b11;
		14'h24f8: color = 2'b11;
		14'h24f9: color = 2'b11;
		14'h24fa: color = 2'b11;
		14'h24fb: color = 2'b11;
		14'h24fc: color = 2'b11;
		14'h24fd: color = 2'b11;
		14'h24fe: color = 2'b11;
		14'h24ff: color = 2'b11;
		14'h2500: color = 2'b11;
		14'h2501: color = 2'b11;
		14'h2502: color = 2'b11;
		14'h2503: color = 2'b11;
		14'h2504: color = 2'b11;
		14'h2505: color = 2'b11;
		14'h2506: color = 2'b11;
		14'h2507: color = 2'b11;
		14'h2508: color = 2'b11;
		14'h2509: color = 2'b11;
		14'h250a: color = 2'b11;
		14'h250b: color = 2'b11;
		14'h250c: color = 2'b11;
		14'h250d: color = 2'b11;
		14'h250e: color = 2'b11;
		14'h250f: color = 2'b11;
		14'h2510: color = 2'b11;
		14'h2511: color = 2'b11;
		14'h2512: color = 2'b11;
		14'h2513: color = 2'b11;
		14'h2514: color = 2'b11;
		14'h2515: color = 2'b11;
		14'h2516: color = 2'b11;
		14'h2517: color = 2'b11;
		14'h2518: color = 2'b11;
		14'h2519: color = 2'b11;
		14'h251a: color = 2'b11;
		14'h251b: color = 2'b11;
		14'h251c: color = 2'b11;
		14'h251d: color = 2'b11;
		14'h251e: color = 2'b11;
		14'h251f: color = 2'b11;
		14'h2520: color = 2'b11;
		14'h2521: color = 2'b11;
		14'h2522: color = 2'b11;
		14'h2523: color = 2'b11;
		14'h2524: color = 2'b11;
		14'h2525: color = 2'b11;
		14'h2526: color = 2'b01;
		14'h2527: color = 2'b00;
		14'h2528: color = 2'b00;
		14'h2529: color = 2'b00;
		14'h252a: color = 2'b10;
		14'h252b: color = 2'b11;
		14'h252c: color = 2'b11;
		14'h252d: color = 2'b10;
		14'h252e: color = 2'b01;
		14'h252f: color = 2'b01;
		14'h2530: color = 2'b01;
		14'h2531: color = 2'b01;
		14'h2532: color = 2'b10;
		14'h2533: color = 2'b01;
		14'h2534: color = 2'b01;
		14'h2535: color = 2'b01;
		14'h2536: color = 2'b01;
		14'h2537: color = 2'b01;
		14'h2538: color = 2'b01;
		14'h2539: color = 2'b10;
		14'h253a: color = 2'b11;
		14'h253b: color = 2'b10;
		14'h253c: color = 2'b01;
		14'h253d: color = 2'b00;
		14'h253e: color = 2'b00;
		14'h253f: color = 2'b00;
		14'h2540: color = 2'b00;
		14'h2541: color = 2'b00;
		14'h2542: color = 2'b00;
		14'h2543: color = 2'b00;
		14'h2544: color = 2'b00;
		14'h2545: color = 2'b01;
		14'h2546: color = 2'b00;
		14'h2547: color = 2'b00;
		14'h2548: color = 2'b00;
		14'h2549: color = 2'b00;
		14'h254a: color = 2'b00;
		14'h254b: color = 2'b00;
		14'h254c: color = 2'b00;
		14'h254d: color = 2'b00;
		14'h254e: color = 2'b00;
		14'h254f: color = 2'b00;
		14'h2550: color = 2'b00;
		14'h2551: color = 2'b00;
		14'h2552: color = 2'b00;
		14'h2553: color = 2'b00;
		14'h2554: color = 2'b00;
		14'h2555: color = 2'b00;
		14'h2556: color = 2'b00;
		14'h2557: color = 2'b00;
		14'h2558: color = 2'b00;
		14'h2559: color = 2'b00;
		14'h255a: color = 2'b01;
		14'h255b: color = 2'b01;
		14'h255c: color = 2'b01;
		14'h255d: color = 2'b00;
		14'h255e: color = 2'b00;
		14'h255f: color = 2'b11;
		14'h2560: color = 2'b11;
		14'h2561: color = 2'b11;
		14'h2562: color = 2'b11;
		14'h2563: color = 2'b11;
		14'h2564: color = 2'b11;
		14'h2565: color = 2'b11;
		14'h2566: color = 2'b11;
		14'h2567: color = 2'b11;
		14'h2568: color = 2'b11;
		14'h2569: color = 2'b11;
		14'h256a: color = 2'b11;
		14'h256b: color = 2'b11;
		14'h256c: color = 2'b11;
		14'h256d: color = 2'b11;
		14'h256e: color = 2'b11;
		14'h256f: color = 2'b11;
		14'h2570: color = 2'b11;
		14'h2571: color = 2'b11;
		14'h2572: color = 2'b11;
		14'h2573: color = 2'b11;
		14'h2574: color = 2'b11;
		14'h2575: color = 2'b11;
		14'h2576: color = 2'b11;
		14'h2577: color = 2'b11;
		14'h2578: color = 2'b11;
		14'h2579: color = 2'b11;
		14'h257a: color = 2'b11;
		14'h257b: color = 2'b11;
		14'h257c: color = 2'b11;
		14'h257d: color = 2'b11;
		14'h257e: color = 2'b11;
		14'h257f: color = 2'b11;
		14'h2580: color = 2'b11;
		14'h2581: color = 2'b11;
		14'h2582: color = 2'b11;
		14'h2583: color = 2'b11;
		14'h2584: color = 2'b11;
		14'h2585: color = 2'b11;
		14'h2586: color = 2'b11;
		14'h2587: color = 2'b11;
		14'h2588: color = 2'b11;
		14'h2589: color = 2'b11;
		14'h258a: color = 2'b11;
		14'h258b: color = 2'b11;
		14'h258c: color = 2'b11;
		14'h258d: color = 2'b11;
		14'h258e: color = 2'b11;
		14'h258f: color = 2'b11;
		14'h2590: color = 2'b11;
		14'h2591: color = 2'b11;
		14'h2592: color = 2'b11;
		14'h2593: color = 2'b11;
		14'h2594: color = 2'b11;
		14'h2595: color = 2'b11;
		14'h2596: color = 2'b11;
		14'h2597: color = 2'b11;
		14'h2598: color = 2'b11;
		14'h2599: color = 2'b11;
		14'h259a: color = 2'b11;
		14'h259b: color = 2'b11;
		14'h259c: color = 2'b11;
		14'h259d: color = 2'b11;
		14'h259e: color = 2'b11;
		14'h259f: color = 2'b11;
		14'h25a0: color = 2'b11;
		14'h25a1: color = 2'b11;
		14'h25a2: color = 2'b11;
		14'h25a3: color = 2'b11;
		14'h25a4: color = 2'b11;
		14'h25a5: color = 2'b01;
		14'h25a6: color = 2'b00;
		14'h25a7: color = 2'b00;
		14'h25a8: color = 2'b00;
		14'h25a9: color = 2'b00;
		14'h25aa: color = 2'b10;
		14'h25ab: color = 2'b10;
		14'h25ac: color = 2'b11;
		14'h25ad: color = 2'b10;
		14'h25ae: color = 2'b10;
		14'h25af: color = 2'b01;
		14'h25b0: color = 2'b10;
		14'h25b1: color = 2'b01;
		14'h25b2: color = 2'b01;
		14'h25b3: color = 2'b01;
		14'h25b4: color = 2'b01;
		14'h25b5: color = 2'b01;
		14'h25b6: color = 2'b01;
		14'h25b7: color = 2'b01;
		14'h25b8: color = 2'b01;
		14'h25b9: color = 2'b10;
		14'h25ba: color = 2'b11;
		14'h25bb: color = 2'b10;
		14'h25bc: color = 2'b01;
		14'h25bd: color = 2'b01;
		14'h25be: color = 2'b00;
		14'h25bf: color = 2'b00;
		14'h25c0: color = 2'b00;
		14'h25c1: color = 2'b00;
		14'h25c2: color = 2'b00;
		14'h25c3: color = 2'b00;
		14'h25c4: color = 2'b00;
		14'h25c5: color = 2'b01;
		14'h25c6: color = 2'b00;
		14'h25c7: color = 2'b00;
		14'h25c8: color = 2'b00;
		14'h25c9: color = 2'b00;
		14'h25ca: color = 2'b00;
		14'h25cb: color = 2'b00;
		14'h25cc: color = 2'b00;
		14'h25cd: color = 2'b00;
		14'h25ce: color = 2'b00;
		14'h25cf: color = 2'b00;
		14'h25d0: color = 2'b00;
		14'h25d1: color = 2'b00;
		14'h25d2: color = 2'b00;
		14'h25d3: color = 2'b00;
		14'h25d4: color = 2'b00;
		14'h25d5: color = 2'b00;
		14'h25d6: color = 2'b00;
		14'h25d7: color = 2'b00;
		14'h25d8: color = 2'b00;
		14'h25d9: color = 2'b00;
		14'h25da: color = 2'b01;
		14'h25db: color = 2'b01;
		14'h25dc: color = 2'b00;
		14'h25dd: color = 2'b00;
		14'h25de: color = 2'b00;
		14'h25df: color = 2'b11;
		14'h25e0: color = 2'b11;
		14'h25e1: color = 2'b11;
		14'h25e2: color = 2'b11;
		14'h25e3: color = 2'b11;
		14'h25e4: color = 2'b11;
		14'h25e5: color = 2'b11;
		14'h25e6: color = 2'b11;
		14'h25e7: color = 2'b11;
		14'h25e8: color = 2'b11;
		14'h25e9: color = 2'b11;
		14'h25ea: color = 2'b11;
		14'h25eb: color = 2'b11;
		14'h25ec: color = 2'b11;
		14'h25ed: color = 2'b11;
		14'h25ee: color = 2'b11;
		14'h25ef: color = 2'b11;
		14'h25f0: color = 2'b11;
		14'h25f1: color = 2'b11;
		14'h25f2: color = 2'b11;
		14'h25f3: color = 2'b11;
		14'h25f4: color = 2'b11;
		14'h25f5: color = 2'b11;
		14'h25f6: color = 2'b11;
		14'h25f7: color = 2'b11;
		14'h25f8: color = 2'b11;
		14'h25f9: color = 2'b11;
		14'h25fa: color = 2'b11;
		14'h25fb: color = 2'b11;
		14'h25fc: color = 2'b11;
		14'h25fd: color = 2'b11;
		14'h25fe: color = 2'b11;
		14'h25ff: color = 2'b11;
		14'h2600: color = 2'b11;
		14'h2601: color = 2'b11;
		14'h2602: color = 2'b11;
		14'h2603: color = 2'b11;
		14'h2604: color = 2'b11;
		14'h2605: color = 2'b11;
		14'h2606: color = 2'b11;
		14'h2607: color = 2'b11;
		14'h2608: color = 2'b11;
		14'h2609: color = 2'b11;
		14'h260a: color = 2'b11;
		14'h260b: color = 2'b11;
		14'h260c: color = 2'b11;
		14'h260d: color = 2'b11;
		14'h260e: color = 2'b11;
		14'h260f: color = 2'b11;
		14'h2610: color = 2'b11;
		14'h2611: color = 2'b11;
		14'h2612: color = 2'b11;
		14'h2613: color = 2'b11;
		14'h2614: color = 2'b11;
		14'h2615: color = 2'b11;
		14'h2616: color = 2'b11;
		14'h2617: color = 2'b11;
		14'h2618: color = 2'b11;
		14'h2619: color = 2'b11;
		14'h261a: color = 2'b11;
		14'h261b: color = 2'b11;
		14'h261c: color = 2'b11;
		14'h261d: color = 2'b11;
		14'h261e: color = 2'b11;
		14'h261f: color = 2'b11;
		14'h2620: color = 2'b11;
		14'h2621: color = 2'b11;
		14'h2622: color = 2'b11;
		14'h2623: color = 2'b11;
		14'h2624: color = 2'b10;
		14'h2625: color = 2'b00;
		14'h2626: color = 2'b01;
		14'h2627: color = 2'b00;
		14'h2628: color = 2'b00;
		14'h2629: color = 2'b00;
		14'h262a: color = 2'b10;
		14'h262b: color = 2'b11;
		14'h262c: color = 2'b11;
		14'h262d: color = 2'b10;
		14'h262e: color = 2'b10;
		14'h262f: color = 2'b00;
		14'h2630: color = 2'b01;
		14'h2631: color = 2'b01;
		14'h2632: color = 2'b01;
		14'h2633: color = 2'b01;
		14'h2634: color = 2'b01;
		14'h2635: color = 2'b01;
		14'h2636: color = 2'b01;
		14'h2637: color = 2'b01;
		14'h2638: color = 2'b01;
		14'h2639: color = 2'b01;
		14'h263a: color = 2'b10;
		14'h263b: color = 2'b01;
		14'h263c: color = 2'b01;
		14'h263d: color = 2'b00;
		14'h263e: color = 2'b00;
		14'h263f: color = 2'b00;
		14'h2640: color = 2'b00;
		14'h2641: color = 2'b00;
		14'h2642: color = 2'b00;
		14'h2643: color = 2'b01;
		14'h2644: color = 2'b01;
		14'h2645: color = 2'b01;
		14'h2646: color = 2'b01;
		14'h2647: color = 2'b01;
		14'h2648: color = 2'b01;
		14'h2649: color = 2'b01;
		14'h264a: color = 2'b01;
		14'h264b: color = 2'b00;
		14'h264c: color = 2'b01;
		14'h264d: color = 2'b01;
		14'h264e: color = 2'b00;
		14'h264f: color = 2'b00;
		14'h2650: color = 2'b00;
		14'h2651: color = 2'b00;
		14'h2652: color = 2'b00;
		14'h2653: color = 2'b00;
		14'h2654: color = 2'b00;
		14'h2655: color = 2'b00;
		14'h2656: color = 2'b00;
		14'h2657: color = 2'b00;
		14'h2658: color = 2'b00;
		14'h2659: color = 2'b00;
		14'h265a: color = 2'b00;
		14'h265b: color = 2'b00;
		14'h265c: color = 2'b00;
		14'h265d: color = 2'b00;
		14'h265e: color = 2'b00;
		14'h265f: color = 2'b11;
		14'h2660: color = 2'b11;
		14'h2661: color = 2'b11;
		14'h2662: color = 2'b11;
		14'h2663: color = 2'b11;
		14'h2664: color = 2'b11;
		14'h2665: color = 2'b11;
		14'h2666: color = 2'b11;
		14'h2667: color = 2'b11;
		14'h2668: color = 2'b11;
		14'h2669: color = 2'b11;
		14'h266a: color = 2'b11;
		14'h266b: color = 2'b11;
		14'h266c: color = 2'b11;
		14'h266d: color = 2'b11;
		14'h266e: color = 2'b11;
		14'h266f: color = 2'b11;
		14'h2670: color = 2'b11;
		14'h2671: color = 2'b11;
		14'h2672: color = 2'b11;
		14'h2673: color = 2'b11;
		14'h2674: color = 2'b11;
		14'h2675: color = 2'b11;
		14'h2676: color = 2'b11;
		14'h2677: color = 2'b11;
		14'h2678: color = 2'b11;
		14'h2679: color = 2'b11;
		14'h267a: color = 2'b11;
		14'h267b: color = 2'b11;
		14'h267c: color = 2'b11;
		14'h267d: color = 2'b11;
		14'h267e: color = 2'b11;
		14'h267f: color = 2'b11;
		14'h2680: color = 2'b11;
		14'h2681: color = 2'b11;
		14'h2682: color = 2'b11;
		14'h2683: color = 2'b11;
		14'h2684: color = 2'b11;
		14'h2685: color = 2'b11;
		14'h2686: color = 2'b11;
		14'h2687: color = 2'b11;
		14'h2688: color = 2'b11;
		14'h2689: color = 2'b11;
		14'h268a: color = 2'b11;
		14'h268b: color = 2'b11;
		14'h268c: color = 2'b11;
		14'h268d: color = 2'b11;
		14'h268e: color = 2'b11;
		14'h268f: color = 2'b11;
		14'h2690: color = 2'b11;
		14'h2691: color = 2'b11;
		14'h2692: color = 2'b11;
		14'h2693: color = 2'b11;
		14'h2694: color = 2'b11;
		14'h2695: color = 2'b11;
		14'h2696: color = 2'b11;
		14'h2697: color = 2'b11;
		14'h2698: color = 2'b11;
		14'h2699: color = 2'b11;
		14'h269a: color = 2'b11;
		14'h269b: color = 2'b11;
		14'h269c: color = 2'b11;
		14'h269d: color = 2'b11;
		14'h269e: color = 2'b11;
		14'h269f: color = 2'b11;
		14'h26a0: color = 2'b11;
		14'h26a1: color = 2'b11;
		14'h26a2: color = 2'b11;
		14'h26a3: color = 2'b11;
		14'h26a4: color = 2'b00;
		14'h26a5: color = 2'b00;
		14'h26a6: color = 2'b00;
		14'h26a7: color = 2'b00;
		14'h26a8: color = 2'b00;
		14'h26a9: color = 2'b00;
		14'h26aa: color = 2'b11;
		14'h26ab: color = 2'b11;
		14'h26ac: color = 2'b11;
		14'h26ad: color = 2'b10;
		14'h26ae: color = 2'b10;
		14'h26af: color = 2'b01;
		14'h26b0: color = 2'b01;
		14'h26b1: color = 2'b01;
		14'h26b2: color = 2'b01;
		14'h26b3: color = 2'b01;
		14'h26b4: color = 2'b01;
		14'h26b5: color = 2'b01;
		14'h26b6: color = 2'b01;
		14'h26b7: color = 2'b00;
		14'h26b8: color = 2'b00;
		14'h26b9: color = 2'b01;
		14'h26ba: color = 2'b10;
		14'h26bb: color = 2'b10;
		14'h26bc: color = 2'b00;
		14'h26bd: color = 2'b00;
		14'h26be: color = 2'b00;
		14'h26bf: color = 2'b00;
		14'h26c0: color = 2'b00;
		14'h26c1: color = 2'b00;
		14'h26c2: color = 2'b01;
		14'h26c3: color = 2'b01;
		14'h26c4: color = 2'b10;
		14'h26c5: color = 2'b10;
		14'h26c6: color = 2'b10;
		14'h26c7: color = 2'b01;
		14'h26c8: color = 2'b01;
		14'h26c9: color = 2'b01;
		14'h26ca: color = 2'b01;
		14'h26cb: color = 2'b01;
		14'h26cc: color = 2'b00;
		14'h26cd: color = 2'b00;
		14'h26ce: color = 2'b00;
		14'h26cf: color = 2'b00;
		14'h26d0: color = 2'b00;
		14'h26d1: color = 2'b00;
		14'h26d2: color = 2'b00;
		14'h26d3: color = 2'b00;
		14'h26d4: color = 2'b00;
		14'h26d5: color = 2'b00;
		14'h26d6: color = 2'b00;
		14'h26d7: color = 2'b00;
		14'h26d8: color = 2'b00;
		14'h26d9: color = 2'b00;
		14'h26da: color = 2'b00;
		14'h26db: color = 2'b00;
		14'h26dc: color = 2'b00;
		14'h26dd: color = 2'b00;
		14'h26de: color = 2'b10;
		14'h26df: color = 2'b11;
		14'h26e0: color = 2'b11;
		14'h26e1: color = 2'b11;
		14'h26e2: color = 2'b11;
		14'h26e3: color = 2'b11;
		14'h26e4: color = 2'b11;
		14'h26e5: color = 2'b11;
		14'h26e6: color = 2'b11;
		14'h26e7: color = 2'b11;
		14'h26e8: color = 2'b11;
		14'h26e9: color = 2'b11;
		14'h26ea: color = 2'b11;
		14'h26eb: color = 2'b11;
		14'h26ec: color = 2'b11;
		14'h26ed: color = 2'b11;
		14'h26ee: color = 2'b11;
		14'h26ef: color = 2'b11;
		14'h26f0: color = 2'b11;
		14'h26f1: color = 2'b11;
		14'h26f2: color = 2'b11;
		14'h26f3: color = 2'b11;
		14'h26f4: color = 2'b11;
		14'h26f5: color = 2'b11;
		14'h26f6: color = 2'b11;
		14'h26f7: color = 2'b11;
		14'h26f8: color = 2'b11;
		14'h26f9: color = 2'b11;
		14'h26fa: color = 2'b11;
		14'h26fb: color = 2'b11;
		14'h26fc: color = 2'b11;
		14'h26fd: color = 2'b11;
		14'h26fe: color = 2'b11;
		14'h26ff: color = 2'b11;
		14'h2700: color = 2'b11;
		14'h2701: color = 2'b11;
		14'h2702: color = 2'b11;
		14'h2703: color = 2'b11;
		14'h2704: color = 2'b11;
		14'h2705: color = 2'b11;
		14'h2706: color = 2'b11;
		14'h2707: color = 2'b11;
		14'h2708: color = 2'b11;
		14'h2709: color = 2'b11;
		14'h270a: color = 2'b11;
		14'h270b: color = 2'b11;
		14'h270c: color = 2'b11;
		14'h270d: color = 2'b11;
		14'h270e: color = 2'b11;
		14'h270f: color = 2'b11;
		14'h2710: color = 2'b11;
		14'h2711: color = 2'b11;
		14'h2712: color = 2'b11;
		14'h2713: color = 2'b11;
		14'h2714: color = 2'b11;
		14'h2715: color = 2'b11;
		14'h2716: color = 2'b11;
		14'h2717: color = 2'b11;
		14'h2718: color = 2'b11;
		14'h2719: color = 2'b11;
		14'h271a: color = 2'b11;
		14'h271b: color = 2'b11;
		14'h271c: color = 2'b11;
		14'h271d: color = 2'b11;
		14'h271e: color = 2'b11;
		14'h271f: color = 2'b11;
		14'h2720: color = 2'b11;
		14'h2721: color = 2'b11;
		14'h2722: color = 2'b11;
		14'h2723: color = 2'b01;
		14'h2724: color = 2'b00;
		14'h2725: color = 2'b01;
		14'h2726: color = 2'b00;
		14'h2727: color = 2'b00;
		14'h2728: color = 2'b00;
		14'h2729: color = 2'b00;
		14'h272a: color = 2'b11;
		14'h272b: color = 2'b11;
		14'h272c: color = 2'b10;
		14'h272d: color = 2'b11;
		14'h272e: color = 2'b10;
		14'h272f: color = 2'b10;
		14'h2730: color = 2'b00;
		14'h2731: color = 2'b01;
		14'h2732: color = 2'b01;
		14'h2733: color = 2'b01;
		14'h2734: color = 2'b01;
		14'h2735: color = 2'b01;
		14'h2736: color = 2'b01;
		14'h2737: color = 2'b00;
		14'h2738: color = 2'b00;
		14'h2739: color = 2'b01;
		14'h273a: color = 2'b01;
		14'h273b: color = 2'b01;
		14'h273c: color = 2'b01;
		14'h273d: color = 2'b00;
		14'h273e: color = 2'b00;
		14'h273f: color = 2'b00;
		14'h2740: color = 2'b00;
		14'h2741: color = 2'b00;
		14'h2742: color = 2'b01;
		14'h2743: color = 2'b10;
		14'h2744: color = 2'b11;
		14'h2745: color = 2'b10;
		14'h2746: color = 2'b10;
		14'h2747: color = 2'b10;
		14'h2748: color = 2'b10;
		14'h2749: color = 2'b10;
		14'h274a: color = 2'b01;
		14'h274b: color = 2'b01;
		14'h274c: color = 2'b01;
		14'h274d: color = 2'b01;
		14'h274e: color = 2'b01;
		14'h274f: color = 2'b01;
		14'h2750: color = 2'b01;
		14'h2751: color = 2'b00;
		14'h2752: color = 2'b00;
		14'h2753: color = 2'b01;
		14'h2754: color = 2'b00;
		14'h2755: color = 2'b00;
		14'h2756: color = 2'b00;
		14'h2757: color = 2'b00;
		14'h2758: color = 2'b00;
		14'h2759: color = 2'b00;
		14'h275a: color = 2'b00;
		14'h275b: color = 2'b00;
		14'h275c: color = 2'b00;
		14'h275d: color = 2'b00;
		14'h275e: color = 2'b11;
		14'h275f: color = 2'b11;
		14'h2760: color = 2'b11;
		14'h2761: color = 2'b11;
		14'h2762: color = 2'b11;
		14'h2763: color = 2'b11;
		14'h2764: color = 2'b11;
		14'h2765: color = 2'b11;
		14'h2766: color = 2'b11;
		14'h2767: color = 2'b11;
		14'h2768: color = 2'b11;
		14'h2769: color = 2'b11;
		14'h276a: color = 2'b11;
		14'h276b: color = 2'b11;
		14'h276c: color = 2'b11;
		14'h276d: color = 2'b11;
		14'h276e: color = 2'b11;
		14'h276f: color = 2'b11;
		14'h2770: color = 2'b11;
		14'h2771: color = 2'b11;
		14'h2772: color = 2'b11;
		14'h2773: color = 2'b11;
		14'h2774: color = 2'b11;
		14'h2775: color = 2'b11;
		14'h2776: color = 2'b11;
		14'h2777: color = 2'b11;
		14'h2778: color = 2'b11;
		14'h2779: color = 2'b11;
		14'h277a: color = 2'b11;
		14'h277b: color = 2'b11;
		14'h277c: color = 2'b11;
		14'h277d: color = 2'b11;
		14'h277e: color = 2'b11;
		14'h277f: color = 2'b11;
		14'h2780: color = 2'b11;
		14'h2781: color = 2'b11;
		14'h2782: color = 2'b11;
		14'h2783: color = 2'b11;
		14'h2784: color = 2'b11;
		14'h2785: color = 2'b11;
		14'h2786: color = 2'b11;
		14'h2787: color = 2'b11;
		14'h2788: color = 2'b11;
		14'h2789: color = 2'b11;
		14'h278a: color = 2'b11;
		14'h278b: color = 2'b11;
		14'h278c: color = 2'b11;
		14'h278d: color = 2'b11;
		14'h278e: color = 2'b11;
		14'h278f: color = 2'b11;
		14'h2790: color = 2'b11;
		14'h2791: color = 2'b11;
		14'h2792: color = 2'b11;
		14'h2793: color = 2'b11;
		14'h2794: color = 2'b11;
		14'h2795: color = 2'b11;
		14'h2796: color = 2'b11;
		14'h2797: color = 2'b11;
		14'h2798: color = 2'b11;
		14'h2799: color = 2'b11;
		14'h279a: color = 2'b11;
		14'h279b: color = 2'b11;
		14'h279c: color = 2'b11;
		14'h279d: color = 2'b11;
		14'h279e: color = 2'b11;
		14'h279f: color = 2'b11;
		14'h27a0: color = 2'b11;
		14'h27a1: color = 2'b11;
		14'h27a2: color = 2'b01;
		14'h27a3: color = 2'b00;
		14'h27a4: color = 2'b00;
		14'h27a5: color = 2'b01;
		14'h27a6: color = 2'b00;
		14'h27a7: color = 2'b00;
		14'h27a8: color = 2'b00;
		14'h27a9: color = 2'b00;
		14'h27aa: color = 2'b11;
		14'h27ab: color = 2'b11;
		14'h27ac: color = 2'b11;
		14'h27ad: color = 2'b10;
		14'h27ae: color = 2'b11;
		14'h27af: color = 2'b10;
		14'h27b0: color = 2'b01;
		14'h27b1: color = 2'b01;
		14'h27b2: color = 2'b01;
		14'h27b3: color = 2'b01;
		14'h27b4: color = 2'b01;
		14'h27b5: color = 2'b00;
		14'h27b6: color = 2'b01;
		14'h27b7: color = 2'b00;
		14'h27b8: color = 2'b00;
		14'h27b9: color = 2'b00;
		14'h27ba: color = 2'b01;
		14'h27bb: color = 2'b01;
		14'h27bc: color = 2'b01;
		14'h27bd: color = 2'b00;
		14'h27be: color = 2'b00;
		14'h27bf: color = 2'b00;
		14'h27c0: color = 2'b00;
		14'h27c1: color = 2'b00;
		14'h27c2: color = 2'b01;
		14'h27c3: color = 2'b10;
		14'h27c4: color = 2'b11;
		14'h27c5: color = 2'b11;
		14'h27c6: color = 2'b11;
		14'h27c7: color = 2'b10;
		14'h27c8: color = 2'b10;
		14'h27c9: color = 2'b10;
		14'h27ca: color = 2'b10;
		14'h27cb: color = 2'b10;
		14'h27cc: color = 2'b10;
		14'h27cd: color = 2'b10;
		14'h27ce: color = 2'b10;
		14'h27cf: color = 2'b01;
		14'h27d0: color = 2'b01;
		14'h27d1: color = 2'b01;
		14'h27d2: color = 2'b01;
		14'h27d3: color = 2'b01;
		14'h27d4: color = 2'b01;
		14'h27d5: color = 2'b00;
		14'h27d6: color = 2'b00;
		14'h27d7: color = 2'b00;
		14'h27d8: color = 2'b00;
		14'h27d9: color = 2'b00;
		14'h27da: color = 2'b00;
		14'h27db: color = 2'b00;
		14'h27dc: color = 2'b00;
		14'h27dd: color = 2'b00;
		14'h27de: color = 2'b11;
		14'h27df: color = 2'b11;
		14'h27e0: color = 2'b11;
		14'h27e1: color = 2'b11;
		14'h27e2: color = 2'b11;
		14'h27e3: color = 2'b11;
		14'h27e4: color = 2'b11;
		14'h27e5: color = 2'b11;
		14'h27e6: color = 2'b11;
		14'h27e7: color = 2'b11;
		14'h27e8: color = 2'b11;
		14'h27e9: color = 2'b11;
		14'h27ea: color = 2'b11;
		14'h27eb: color = 2'b11;
		14'h27ec: color = 2'b11;
		14'h27ed: color = 2'b11;
		14'h27ee: color = 2'b11;
		14'h27ef: color = 2'b11;
		14'h27f0: color = 2'b11;
		14'h27f1: color = 2'b11;
		14'h27f2: color = 2'b11;
		14'h27f3: color = 2'b11;
		14'h27f4: color = 2'b11;
		14'h27f5: color = 2'b11;
		14'h27f6: color = 2'b11;
		14'h27f7: color = 2'b11;
		14'h27f8: color = 2'b11;
		14'h27f9: color = 2'b11;
		14'h27fa: color = 2'b11;
		14'h27fb: color = 2'b11;
		14'h27fc: color = 2'b11;
		14'h27fd: color = 2'b11;
		14'h27fe: color = 2'b11;
		14'h27ff: color = 2'b11;
		14'h2800: color = 2'b11;
		14'h2801: color = 2'b11;
		14'h2802: color = 2'b11;
		14'h2803: color = 2'b11;
		14'h2804: color = 2'b11;
		14'h2805: color = 2'b11;
		14'h2806: color = 2'b11;
		14'h2807: color = 2'b11;
		14'h2808: color = 2'b11;
		14'h2809: color = 2'b11;
		14'h280a: color = 2'b11;
		14'h280b: color = 2'b11;
		14'h280c: color = 2'b11;
		14'h280d: color = 2'b11;
		14'h280e: color = 2'b11;
		14'h280f: color = 2'b11;
		14'h2810: color = 2'b11;
		14'h2811: color = 2'b11;
		14'h2812: color = 2'b11;
		14'h2813: color = 2'b11;
		14'h2814: color = 2'b11;
		14'h2815: color = 2'b11;
		14'h2816: color = 2'b11;
		14'h2817: color = 2'b11;
		14'h2818: color = 2'b11;
		14'h2819: color = 2'b11;
		14'h281a: color = 2'b11;
		14'h281b: color = 2'b11;
		14'h281c: color = 2'b11;
		14'h281d: color = 2'b11;
		14'h281e: color = 2'b11;
		14'h281f: color = 2'b11;
		14'h2820: color = 2'b11;
		14'h2821: color = 2'b00;
		14'h2822: color = 2'b01;
		14'h2823: color = 2'b00;
		14'h2824: color = 2'b01;
		14'h2825: color = 2'b00;
		14'h2826: color = 2'b00;
		14'h2827: color = 2'b01;
		14'h2828: color = 2'b01;
		14'h2829: color = 2'b00;
		14'h282a: color = 2'b11;
		14'h282b: color = 2'b11;
		14'h282c: color = 2'b11;
		14'h282d: color = 2'b11;
		14'h282e: color = 2'b10;
		14'h282f: color = 2'b11;
		14'h2830: color = 2'b10;
		14'h2831: color = 2'b01;
		14'h2832: color = 2'b01;
		14'h2833: color = 2'b00;
		14'h2834: color = 2'b01;
		14'h2835: color = 2'b01;
		14'h2836: color = 2'b00;
		14'h2837: color = 2'b00;
		14'h2838: color = 2'b00;
		14'h2839: color = 2'b01;
		14'h283a: color = 2'b01;
		14'h283b: color = 2'b01;
		14'h283c: color = 2'b00;
		14'h283d: color = 2'b01;
		14'h283e: color = 2'b01;
		14'h283f: color = 2'b00;
		14'h2840: color = 2'b00;
		14'h2841: color = 2'b01;
		14'h2842: color = 2'b01;
		14'h2843: color = 2'b01;
		14'h2844: color = 2'b10;
		14'h2845: color = 2'b10;
		14'h2846: color = 2'b10;
		14'h2847: color = 2'b10;
		14'h2848: color = 2'b10;
		14'h2849: color = 2'b10;
		14'h284a: color = 2'b10;
		14'h284b: color = 2'b01;
		14'h284c: color = 2'b10;
		14'h284d: color = 2'b01;
		14'h284e: color = 2'b01;
		14'h284f: color = 2'b01;
		14'h2850: color = 2'b01;
		14'h2851: color = 2'b01;
		14'h2852: color = 2'b01;
		14'h2853: color = 2'b01;
		14'h2854: color = 2'b00;
		14'h2855: color = 2'b00;
		14'h2856: color = 2'b00;
		14'h2857: color = 2'b00;
		14'h2858: color = 2'b00;
		14'h2859: color = 2'b00;
		14'h285a: color = 2'b00;
		14'h285b: color = 2'b00;
		14'h285c: color = 2'b00;
		14'h285d: color = 2'b10;
		14'h285e: color = 2'b11;
		14'h285f: color = 2'b11;
		14'h2860: color = 2'b11;
		14'h2861: color = 2'b11;
		14'h2862: color = 2'b11;
		14'h2863: color = 2'b11;
		14'h2864: color = 2'b11;
		14'h2865: color = 2'b11;
		14'h2866: color = 2'b11;
		14'h2867: color = 2'b11;
		14'h2868: color = 2'b11;
		14'h2869: color = 2'b11;
		14'h286a: color = 2'b11;
		14'h286b: color = 2'b11;
		14'h286c: color = 2'b11;
		14'h286d: color = 2'b11;
		14'h286e: color = 2'b11;
		14'h286f: color = 2'b11;
		14'h2870: color = 2'b11;
		14'h2871: color = 2'b11;
		14'h2872: color = 2'b11;
		14'h2873: color = 2'b11;
		14'h2874: color = 2'b11;
		14'h2875: color = 2'b11;
		14'h2876: color = 2'b11;
		14'h2877: color = 2'b11;
		14'h2878: color = 2'b11;
		14'h2879: color = 2'b11;
		14'h287a: color = 2'b11;
		14'h287b: color = 2'b11;
		14'h287c: color = 2'b11;
		14'h287d: color = 2'b11;
		14'h287e: color = 2'b11;
		14'h287f: color = 2'b11;
		14'h2880: color = 2'b11;
		14'h2881: color = 2'b11;
		14'h2882: color = 2'b11;
		14'h2883: color = 2'b11;
		14'h2884: color = 2'b11;
		14'h2885: color = 2'b11;
		14'h2886: color = 2'b11;
		14'h2887: color = 2'b11;
		14'h2888: color = 2'b11;
		14'h2889: color = 2'b11;
		14'h288a: color = 2'b11;
		14'h288b: color = 2'b11;
		14'h288c: color = 2'b11;
		14'h288d: color = 2'b11;
		14'h288e: color = 2'b11;
		14'h288f: color = 2'b11;
		14'h2890: color = 2'b11;
		14'h2891: color = 2'b11;
		14'h2892: color = 2'b11;
		14'h2893: color = 2'b11;
		14'h2894: color = 2'b11;
		14'h2895: color = 2'b11;
		14'h2896: color = 2'b11;
		14'h2897: color = 2'b11;
		14'h2898: color = 2'b11;
		14'h2899: color = 2'b11;
		14'h289a: color = 2'b11;
		14'h289b: color = 2'b11;
		14'h289c: color = 2'b11;
		14'h289d: color = 2'b11;
		14'h289e: color = 2'b11;
		14'h289f: color = 2'b01;
		14'h28a0: color = 2'b00;
		14'h28a1: color = 2'b00;
		14'h28a2: color = 2'b00;
		14'h28a3: color = 2'b00;
		14'h28a4: color = 2'b01;
		14'h28a5: color = 2'b01;
		14'h28a6: color = 2'b00;
		14'h28a7: color = 2'b00;
		14'h28a8: color = 2'b00;
		14'h28a9: color = 2'b00;
		14'h28aa: color = 2'b11;
		14'h28ab: color = 2'b11;
		14'h28ac: color = 2'b11;
		14'h28ad: color = 2'b11;
		14'h28ae: color = 2'b10;
		14'h28af: color = 2'b11;
		14'h28b0: color = 2'b10;
		14'h28b1: color = 2'b01;
		14'h28b2: color = 2'b00;
		14'h28b3: color = 2'b01;
		14'h28b4: color = 2'b00;
		14'h28b5: color = 2'b01;
		14'h28b6: color = 2'b01;
		14'h28b7: color = 2'b00;
		14'h28b8: color = 2'b00;
		14'h28b9: color = 2'b00;
		14'h28ba: color = 2'b00;
		14'h28bb: color = 2'b01;
		14'h28bc: color = 2'b01;
		14'h28bd: color = 2'b00;
		14'h28be: color = 2'b00;
		14'h28bf: color = 2'b01;
		14'h28c0: color = 2'b00;
		14'h28c1: color = 2'b00;
		14'h28c2: color = 2'b01;
		14'h28c3: color = 2'b01;
		14'h28c4: color = 2'b01;
		14'h28c5: color = 2'b01;
		14'h28c6: color = 2'b01;
		14'h28c7: color = 2'b01;
		14'h28c8: color = 2'b01;
		14'h28c9: color = 2'b01;
		14'h28ca: color = 2'b01;
		14'h28cb: color = 2'b00;
		14'h28cc: color = 2'b00;
		14'h28cd: color = 2'b00;
		14'h28ce: color = 2'b01;
		14'h28cf: color = 2'b01;
		14'h28d0: color = 2'b00;
		14'h28d1: color = 2'b01;
		14'h28d2: color = 2'b01;
		14'h28d3: color = 2'b01;
		14'h28d4: color = 2'b00;
		14'h28d5: color = 2'b00;
		14'h28d6: color = 2'b00;
		14'h28d7: color = 2'b00;
		14'h28d8: color = 2'b00;
		14'h28d9: color = 2'b00;
		14'h28da: color = 2'b00;
		14'h28db: color = 2'b00;
		14'h28dc: color = 2'b00;
		14'h28dd: color = 2'b11;
		14'h28de: color = 2'b11;
		14'h28df: color = 2'b11;
		14'h28e0: color = 2'b11;
		14'h28e1: color = 2'b11;
		14'h28e2: color = 2'b11;
		14'h28e3: color = 2'b11;
		14'h28e4: color = 2'b11;
		14'h28e5: color = 2'b11;
		14'h28e6: color = 2'b11;
		14'h28e7: color = 2'b11;
		14'h28e8: color = 2'b11;
		14'h28e9: color = 2'b11;
		14'h28ea: color = 2'b11;
		14'h28eb: color = 2'b11;
		14'h28ec: color = 2'b11;
		14'h28ed: color = 2'b11;
		14'h28ee: color = 2'b11;
		14'h28ef: color = 2'b11;
		14'h28f0: color = 2'b11;
		14'h28f1: color = 2'b11;
		14'h28f2: color = 2'b11;
		14'h28f3: color = 2'b11;
		14'h28f4: color = 2'b11;
		14'h28f5: color = 2'b11;
		14'h28f6: color = 2'b11;
		14'h28f7: color = 2'b11;
		14'h28f8: color = 2'b11;
		14'h28f9: color = 2'b11;
		14'h28fa: color = 2'b11;
		14'h28fb: color = 2'b11;
		14'h28fc: color = 2'b11;
		14'h28fd: color = 2'b11;
		14'h28fe: color = 2'b11;
		14'h28ff: color = 2'b11;
		14'h2900: color = 2'b11;
		14'h2901: color = 2'b11;
		14'h2902: color = 2'b11;
		14'h2903: color = 2'b11;
		14'h2904: color = 2'b11;
		14'h2905: color = 2'b11;
		14'h2906: color = 2'b11;
		14'h2907: color = 2'b11;
		14'h2908: color = 2'b11;
		14'h2909: color = 2'b11;
		14'h290a: color = 2'b11;
		14'h290b: color = 2'b11;
		14'h290c: color = 2'b11;
		14'h290d: color = 2'b11;
		14'h290e: color = 2'b11;
		14'h290f: color = 2'b11;
		14'h2910: color = 2'b11;
		14'h2911: color = 2'b11;
		14'h2912: color = 2'b11;
		14'h2913: color = 2'b11;
		14'h2914: color = 2'b11;
		14'h2915: color = 2'b11;
		14'h2916: color = 2'b11;
		14'h2917: color = 2'b11;
		14'h2918: color = 2'b11;
		14'h2919: color = 2'b11;
		14'h291a: color = 2'b11;
		14'h291b: color = 2'b11;
		14'h291c: color = 2'b11;
		14'h291d: color = 2'b11;
		14'h291e: color = 2'b01;
		14'h291f: color = 2'b00;
		14'h2920: color = 2'b00;
		14'h2921: color = 2'b01;
		14'h2922: color = 2'b01;
		14'h2923: color = 2'b00;
		14'h2924: color = 2'b00;
		14'h2925: color = 2'b00;
		14'h2926: color = 2'b00;
		14'h2927: color = 2'b00;
		14'h2928: color = 2'b00;
		14'h2929: color = 2'b00;
		14'h292a: color = 2'b10;
		14'h292b: color = 2'b11;
		14'h292c: color = 2'b11;
		14'h292d: color = 2'b11;
		14'h292e: color = 2'b11;
		14'h292f: color = 2'b10;
		14'h2930: color = 2'b10;
		14'h2931: color = 2'b10;
		14'h2932: color = 2'b01;
		14'h2933: color = 2'b00;
		14'h2934: color = 2'b01;
		14'h2935: color = 2'b00;
		14'h2936: color = 2'b01;
		14'h2937: color = 2'b00;
		14'h2938: color = 2'b00;
		14'h2939: color = 2'b00;
		14'h293a: color = 2'b00;
		14'h293b: color = 2'b00;
		14'h293c: color = 2'b00;
		14'h293d: color = 2'b01;
		14'h293e: color = 2'b00;
		14'h293f: color = 2'b01;
		14'h2940: color = 2'b00;
		14'h2941: color = 2'b00;
		14'h2942: color = 2'b01;
		14'h2943: color = 2'b00;
		14'h2944: color = 2'b01;
		14'h2945: color = 2'b01;
		14'h2946: color = 2'b00;
		14'h2947: color = 2'b01;
		14'h2948: color = 2'b01;
		14'h2949: color = 2'b00;
		14'h294a: color = 2'b00;
		14'h294b: color = 2'b00;
		14'h294c: color = 2'b00;
		14'h294d: color = 2'b00;
		14'h294e: color = 2'b01;
		14'h294f: color = 2'b00;
		14'h2950: color = 2'b00;
		14'h2951: color = 2'b00;
		14'h2952: color = 2'b00;
		14'h2953: color = 2'b00;
		14'h2954: color = 2'b00;
		14'h2955: color = 2'b00;
		14'h2956: color = 2'b00;
		14'h2957: color = 2'b00;
		14'h2958: color = 2'b00;
		14'h2959: color = 2'b00;
		14'h295a: color = 2'b00;
		14'h295b: color = 2'b00;
		14'h295c: color = 2'b10;
		14'h295d: color = 2'b11;
		14'h295e: color = 2'b11;
		14'h295f: color = 2'b11;
		14'h2960: color = 2'b11;
		14'h2961: color = 2'b11;
		14'h2962: color = 2'b11;
		14'h2963: color = 2'b11;
		14'h2964: color = 2'b11;
		14'h2965: color = 2'b11;
		14'h2966: color = 2'b11;
		14'h2967: color = 2'b11;
		14'h2968: color = 2'b11;
		14'h2969: color = 2'b11;
		14'h296a: color = 2'b11;
		14'h296b: color = 2'b11;
		14'h296c: color = 2'b11;
		14'h296d: color = 2'b11;
		14'h296e: color = 2'b11;
		14'h296f: color = 2'b11;
		14'h2970: color = 2'b11;
		14'h2971: color = 2'b11;
		14'h2972: color = 2'b11;
		14'h2973: color = 2'b11;
		14'h2974: color = 2'b11;
		14'h2975: color = 2'b11;
		14'h2976: color = 2'b11;
		14'h2977: color = 2'b11;
		14'h2978: color = 2'b11;
		14'h2979: color = 2'b11;
		14'h297a: color = 2'b11;
		14'h297b: color = 2'b11;
		14'h297c: color = 2'b11;
		14'h297d: color = 2'b11;
		14'h297e: color = 2'b11;
		14'h297f: color = 2'b11;
		14'h2980: color = 2'b11;
		14'h2981: color = 2'b11;
		14'h2982: color = 2'b11;
		14'h2983: color = 2'b11;
		14'h2984: color = 2'b11;
		14'h2985: color = 2'b11;
		14'h2986: color = 2'b11;
		14'h2987: color = 2'b11;
		14'h2988: color = 2'b11;
		14'h2989: color = 2'b11;
		14'h298a: color = 2'b11;
		14'h298b: color = 2'b11;
		14'h298c: color = 2'b11;
		14'h298d: color = 2'b11;
		14'h298e: color = 2'b11;
		14'h298f: color = 2'b11;
		14'h2990: color = 2'b11;
		14'h2991: color = 2'b11;
		14'h2992: color = 2'b11;
		14'h2993: color = 2'b11;
		14'h2994: color = 2'b11;
		14'h2995: color = 2'b11;
		14'h2996: color = 2'b11;
		14'h2997: color = 2'b11;
		14'h2998: color = 2'b11;
		14'h2999: color = 2'b11;
		14'h299a: color = 2'b11;
		14'h299b: color = 2'b11;
		14'h299c: color = 2'b10;
		14'h299d: color = 2'b01;
		14'h299e: color = 2'b00;
		14'h299f: color = 2'b01;
		14'h29a0: color = 2'b00;
		14'h29a1: color = 2'b00;
		14'h29a2: color = 2'b00;
		14'h29a3: color = 2'b01;
		14'h29a4: color = 2'b00;
		14'h29a5: color = 2'b01;
		14'h29a6: color = 2'b01;
		14'h29a7: color = 2'b00;
		14'h29a8: color = 2'b00;
		14'h29a9: color = 2'b00;
		14'h29aa: color = 2'b01;
		14'h29ab: color = 2'b11;
		14'h29ac: color = 2'b11;
		14'h29ad: color = 2'b11;
		14'h29ae: color = 2'b11;
		14'h29af: color = 2'b10;
		14'h29b0: color = 2'b11;
		14'h29b1: color = 2'b11;
		14'h29b2: color = 2'b10;
		14'h29b3: color = 2'b00;
		14'h29b4: color = 2'b00;
		14'h29b5: color = 2'b00;
		14'h29b6: color = 2'b00;
		14'h29b7: color = 2'b00;
		14'h29b8: color = 2'b00;
		14'h29b9: color = 2'b00;
		14'h29ba: color = 2'b01;
		14'h29bb: color = 2'b00;
		14'h29bc: color = 2'b01;
		14'h29bd: color = 2'b00;
		14'h29be: color = 2'b00;
		14'h29bf: color = 2'b00;
		14'h29c0: color = 2'b00;
		14'h29c1: color = 2'b00;
		14'h29c2: color = 2'b00;
		14'h29c3: color = 2'b00;
		14'h29c4: color = 2'b00;
		14'h29c5: color = 2'b01;
		14'h29c6: color = 2'b00;
		14'h29c7: color = 2'b00;
		14'h29c8: color = 2'b00;
		14'h29c9: color = 2'b00;
		14'h29ca: color = 2'b00;
		14'h29cb: color = 2'b00;
		14'h29cc: color = 2'b00;
		14'h29cd: color = 2'b00;
		14'h29ce: color = 2'b00;
		14'h29cf: color = 2'b00;
		14'h29d0: color = 2'b01;
		14'h29d1: color = 2'b00;
		14'h29d2: color = 2'b00;
		14'h29d3: color = 2'b00;
		14'h29d4: color = 2'b00;
		14'h29d5: color = 2'b00;
		14'h29d6: color = 2'b00;
		14'h29d7: color = 2'b00;
		14'h29d8: color = 2'b00;
		14'h29d9: color = 2'b00;
		14'h29da: color = 2'b00;
		14'h29db: color = 2'b00;
		14'h29dc: color = 2'b11;
		14'h29dd: color = 2'b11;
		14'h29de: color = 2'b11;
		14'h29df: color = 2'b11;
		14'h29e0: color = 2'b11;
		14'h29e1: color = 2'b11;
		14'h29e2: color = 2'b11;
		14'h29e3: color = 2'b11;
		14'h29e4: color = 2'b11;
		14'h29e5: color = 2'b11;
		14'h29e6: color = 2'b11;
		14'h29e7: color = 2'b11;
		14'h29e8: color = 2'b11;
		14'h29e9: color = 2'b11;
		14'h29ea: color = 2'b11;
		14'h29eb: color = 2'b11;
		14'h29ec: color = 2'b11;
		14'h29ed: color = 2'b11;
		14'h29ee: color = 2'b11;
		14'h29ef: color = 2'b11;
		14'h29f0: color = 2'b11;
		14'h29f1: color = 2'b11;
		14'h29f2: color = 2'b11;
		14'h29f3: color = 2'b11;
		14'h29f4: color = 2'b11;
		14'h29f5: color = 2'b11;
		14'h29f6: color = 2'b11;
		14'h29f7: color = 2'b11;
		14'h29f8: color = 2'b11;
		14'h29f9: color = 2'b11;
		14'h29fa: color = 2'b11;
		14'h29fb: color = 2'b11;
		14'h29fc: color = 2'b11;
		14'h29fd: color = 2'b11;
		14'h29fe: color = 2'b11;
		14'h29ff: color = 2'b11;
		14'h2a00: color = 2'b11;
		14'h2a01: color = 2'b11;
		14'h2a02: color = 2'b11;
		14'h2a03: color = 2'b11;
		14'h2a04: color = 2'b11;
		14'h2a05: color = 2'b11;
		14'h2a06: color = 2'b11;
		14'h2a07: color = 2'b11;
		14'h2a08: color = 2'b11;
		14'h2a09: color = 2'b11;
		14'h2a0a: color = 2'b11;
		14'h2a0b: color = 2'b11;
		14'h2a0c: color = 2'b11;
		14'h2a0d: color = 2'b11;
		14'h2a0e: color = 2'b11;
		14'h2a0f: color = 2'b11;
		14'h2a10: color = 2'b11;
		14'h2a11: color = 2'b11;
		14'h2a12: color = 2'b11;
		14'h2a13: color = 2'b11;
		14'h2a14: color = 2'b11;
		14'h2a15: color = 2'b11;
		14'h2a16: color = 2'b11;
		14'h2a17: color = 2'b11;
		14'h2a18: color = 2'b11;
		14'h2a19: color = 2'b11;
		14'h2a1a: color = 2'b11;
		14'h2a1b: color = 2'b10;
		14'h2a1c: color = 2'b01;
		14'h2a1d: color = 2'b00;
		14'h2a1e: color = 2'b00;
		14'h2a1f: color = 2'b00;
		14'h2a20: color = 2'b00;
		14'h2a21: color = 2'b00;
		14'h2a22: color = 2'b00;
		14'h2a23: color = 2'b00;
		14'h2a24: color = 2'b00;
		14'h2a25: color = 2'b01;
		14'h2a26: color = 2'b00;
		14'h2a27: color = 2'b01;
		14'h2a28: color = 2'b01;
		14'h2a29: color = 2'b00;
		14'h2a2a: color = 2'b00;
		14'h2a2b: color = 2'b11;
		14'h2a2c: color = 2'b11;
		14'h2a2d: color = 2'b11;
		14'h2a2e: color = 2'b11;
		14'h2a2f: color = 2'b11;
		14'h2a30: color = 2'b10;
		14'h2a31: color = 2'b10;
		14'h2a32: color = 2'b10;
		14'h2a33: color = 2'b01;
		14'h2a34: color = 2'b00;
		14'h2a35: color = 2'b00;
		14'h2a36: color = 2'b01;
		14'h2a37: color = 2'b00;
		14'h2a38: color = 2'b00;
		14'h2a39: color = 2'b00;
		14'h2a3a: color = 2'b00;
		14'h2a3b: color = 2'b01;
		14'h2a3c: color = 2'b00;
		14'h2a3d: color = 2'b00;
		14'h2a3e: color = 2'b01;
		14'h2a3f: color = 2'b00;
		14'h2a40: color = 2'b00;
		14'h2a41: color = 2'b01;
		14'h2a42: color = 2'b00;
		14'h2a43: color = 2'b00;
		14'h2a44: color = 2'b00;
		14'h2a45: color = 2'b00;
		14'h2a46: color = 2'b00;
		14'h2a47: color = 2'b00;
		14'h2a48: color = 2'b00;
		14'h2a49: color = 2'b00;
		14'h2a4a: color = 2'b00;
		14'h2a4b: color = 2'b00;
		14'h2a4c: color = 2'b00;
		14'h2a4d: color = 2'b00;
		14'h2a4e: color = 2'b00;
		14'h2a4f: color = 2'b01;
		14'h2a50: color = 2'b00;
		14'h2a51: color = 2'b00;
		14'h2a52: color = 2'b00;
		14'h2a53: color = 2'b00;
		14'h2a54: color = 2'b00;
		14'h2a55: color = 2'b00;
		14'h2a56: color = 2'b00;
		14'h2a57: color = 2'b00;
		14'h2a58: color = 2'b00;
		14'h2a59: color = 2'b00;
		14'h2a5a: color = 2'b00;
		14'h2a5b: color = 2'b10;
		14'h2a5c: color = 2'b11;
		14'h2a5d: color = 2'b11;
		14'h2a5e: color = 2'b11;
		14'h2a5f: color = 2'b11;
		14'h2a60: color = 2'b11;
		14'h2a61: color = 2'b11;
		14'h2a62: color = 2'b11;
		14'h2a63: color = 2'b11;
		14'h2a64: color = 2'b11;
		14'h2a65: color = 2'b11;
		14'h2a66: color = 2'b11;
		14'h2a67: color = 2'b11;
		14'h2a68: color = 2'b11;
		14'h2a69: color = 2'b11;
		14'h2a6a: color = 2'b11;
		14'h2a6b: color = 2'b11;
		14'h2a6c: color = 2'b11;
		14'h2a6d: color = 2'b11;
		14'h2a6e: color = 2'b11;
		14'h2a6f: color = 2'b11;
		14'h2a70: color = 2'b11;
		14'h2a71: color = 2'b11;
		14'h2a72: color = 2'b11;
		14'h2a73: color = 2'b11;
		14'h2a74: color = 2'b11;
		14'h2a75: color = 2'b11;
		14'h2a76: color = 2'b11;
		14'h2a77: color = 2'b11;
		14'h2a78: color = 2'b11;
		14'h2a79: color = 2'b11;
		14'h2a7a: color = 2'b11;
		14'h2a7b: color = 2'b11;
		14'h2a7c: color = 2'b11;
		14'h2a7d: color = 2'b11;
		14'h2a7e: color = 2'b11;
		14'h2a7f: color = 2'b11;
		14'h2a80: color = 2'b11;
		14'h2a81: color = 2'b11;
		14'h2a82: color = 2'b11;
		14'h2a83: color = 2'b11;
		14'h2a84: color = 2'b11;
		14'h2a85: color = 2'b11;
		14'h2a86: color = 2'b11;
		14'h2a87: color = 2'b11;
		14'h2a88: color = 2'b11;
		14'h2a89: color = 2'b11;
		14'h2a8a: color = 2'b11;
		14'h2a8b: color = 2'b11;
		14'h2a8c: color = 2'b11;
		14'h2a8d: color = 2'b11;
		14'h2a8e: color = 2'b11;
		14'h2a8f: color = 2'b11;
		14'h2a90: color = 2'b11;
		14'h2a91: color = 2'b11;
		14'h2a92: color = 2'b11;
		14'h2a93: color = 2'b11;
		14'h2a94: color = 2'b11;
		14'h2a95: color = 2'b11;
		14'h2a96: color = 2'b11;
		14'h2a97: color = 2'b11;
		14'h2a98: color = 2'b11;
		14'h2a99: color = 2'b10;
		14'h2a9a: color = 2'b01;
		14'h2a9b: color = 2'b00;
		14'h2a9c: color = 2'b00;
		14'h2a9d: color = 2'b00;
		14'h2a9e: color = 2'b00;
		14'h2a9f: color = 2'b00;
		14'h2aa0: color = 2'b00;
		14'h2aa1: color = 2'b00;
		14'h2aa2: color = 2'b01;
		14'h2aa3: color = 2'b00;
		14'h2aa4: color = 2'b01;
		14'h2aa5: color = 2'b00;
		14'h2aa6: color = 2'b00;
		14'h2aa7: color = 2'b00;
		14'h2aa8: color = 2'b00;
		14'h2aa9: color = 2'b00;
		14'h2aaa: color = 2'b00;
		14'h2aab: color = 2'b10;
		14'h2aac: color = 2'b11;
		14'h2aad: color = 2'b11;
		14'h2aae: color = 2'b11;
		14'h2aaf: color = 2'b11;
		14'h2ab0: color = 2'b11;
		14'h2ab1: color = 2'b10;
		14'h2ab2: color = 2'b10;
		14'h2ab3: color = 2'b10;
		14'h2ab4: color = 2'b01;
		14'h2ab5: color = 2'b00;
		14'h2ab6: color = 2'b00;
		14'h2ab7: color = 2'b00;
		14'h2ab8: color = 2'b00;
		14'h2ab9: color = 2'b00;
		14'h2aba: color = 2'b00;
		14'h2abb: color = 2'b00;
		14'h2abc: color = 2'b00;
		14'h2abd: color = 2'b00;
		14'h2abe: color = 2'b00;
		14'h2abf: color = 2'b00;
		14'h2ac0: color = 2'b00;
		14'h2ac1: color = 2'b00;
		14'h2ac2: color = 2'b00;
		14'h2ac3: color = 2'b00;
		14'h2ac4: color = 2'b00;
		14'h2ac5: color = 2'b00;
		14'h2ac6: color = 2'b00;
		14'h2ac7: color = 2'b00;
		14'h2ac8: color = 2'b00;
		14'h2ac9: color = 2'b00;
		14'h2aca: color = 2'b00;
		14'h2acb: color = 2'b00;
		14'h2acc: color = 2'b00;
		14'h2acd: color = 2'b00;
		14'h2ace: color = 2'b00;
		14'h2acf: color = 2'b00;
		14'h2ad0: color = 2'b00;
		14'h2ad1: color = 2'b00;
		14'h2ad2: color = 2'b00;
		14'h2ad3: color = 2'b00;
		14'h2ad4: color = 2'b00;
		14'h2ad5: color = 2'b00;
		14'h2ad6: color = 2'b00;
		14'h2ad7: color = 2'b00;
		14'h2ad8: color = 2'b00;
		14'h2ad9: color = 2'b00;
		14'h2ada: color = 2'b10;
		14'h2adb: color = 2'b11;
		14'h2adc: color = 2'b11;
		14'h2add: color = 2'b11;
		14'h2ade: color = 2'b11;
		14'h2adf: color = 2'b11;
		14'h2ae0: color = 2'b11;
		14'h2ae1: color = 2'b11;
		14'h2ae2: color = 2'b11;
		14'h2ae3: color = 2'b11;
		14'h2ae4: color = 2'b11;
		14'h2ae5: color = 2'b11;
		14'h2ae6: color = 2'b11;
		14'h2ae7: color = 2'b11;
		14'h2ae8: color = 2'b11;
		14'h2ae9: color = 2'b11;
		14'h2aea: color = 2'b11;
		14'h2aeb: color = 2'b11;
		14'h2aec: color = 2'b11;
		14'h2aed: color = 2'b11;
		14'h2aee: color = 2'b11;
		14'h2aef: color = 2'b11;
		14'h2af0: color = 2'b11;
		14'h2af1: color = 2'b11;
		14'h2af2: color = 2'b11;
		14'h2af3: color = 2'b11;
		14'h2af4: color = 2'b11;
		14'h2af5: color = 2'b11;
		14'h2af6: color = 2'b11;
		14'h2af7: color = 2'b11;
		14'h2af8: color = 2'b11;
		14'h2af9: color = 2'b11;
		14'h2afa: color = 2'b11;
		14'h2afb: color = 2'b11;
		14'h2afc: color = 2'b11;
		14'h2afd: color = 2'b11;
		14'h2afe: color = 2'b11;
		14'h2aff: color = 2'b11;
		14'h2b00: color = 2'b11;
		14'h2b01: color = 2'b11;
		14'h2b02: color = 2'b11;
		14'h2b03: color = 2'b11;
		14'h2b04: color = 2'b11;
		14'h2b05: color = 2'b11;
		14'h2b06: color = 2'b11;
		14'h2b07: color = 2'b11;
		14'h2b08: color = 2'b11;
		14'h2b09: color = 2'b11;
		14'h2b0a: color = 2'b11;
		14'h2b0b: color = 2'b11;
		14'h2b0c: color = 2'b11;
		14'h2b0d: color = 2'b11;
		14'h2b0e: color = 2'b11;
		14'h2b0f: color = 2'b11;
		14'h2b10: color = 2'b11;
		14'h2b11: color = 2'b11;
		14'h2b12: color = 2'b11;
		14'h2b13: color = 2'b11;
		14'h2b14: color = 2'b11;
		14'h2b15: color = 2'b11;
		14'h2b16: color = 2'b10;
		14'h2b17: color = 2'b01;
		14'h2b18: color = 2'b01;
		14'h2b19: color = 2'b00;
		14'h2b1a: color = 2'b00;
		14'h2b1b: color = 2'b00;
		14'h2b1c: color = 2'b01;
		14'h2b1d: color = 2'b00;
		14'h2b1e: color = 2'b00;
		14'h2b1f: color = 2'b00;
		14'h2b20: color = 2'b00;
		14'h2b21: color = 2'b00;
		14'h2b22: color = 2'b00;
		14'h2b23: color = 2'b00;
		14'h2b24: color = 2'b00;
		14'h2b25: color = 2'b01;
		14'h2b26: color = 2'b00;
		14'h2b27: color = 2'b01;
		14'h2b28: color = 2'b01;
		14'h2b29: color = 2'b00;
		14'h2b2a: color = 2'b00;
		14'h2b2b: color = 2'b01;
		14'h2b2c: color = 2'b11;
		14'h2b2d: color = 2'b11;
		14'h2b2e: color = 2'b11;
		14'h2b2f: color = 2'b11;
		14'h2b30: color = 2'b11;
		14'h2b31: color = 2'b10;
		14'h2b32: color = 2'b10;
		14'h2b33: color = 2'b10;
		14'h2b34: color = 2'b01;
		14'h2b35: color = 2'b01;
		14'h2b36: color = 2'b00;
		14'h2b37: color = 2'b00;
		14'h2b38: color = 2'b00;
		14'h2b39: color = 2'b00;
		14'h2b3a: color = 2'b00;
		14'h2b3b: color = 2'b00;
		14'h2b3c: color = 2'b00;
		14'h2b3d: color = 2'b00;
		14'h2b3e: color = 2'b00;
		14'h2b3f: color = 2'b01;
		14'h2b40: color = 2'b00;
		14'h2b41: color = 2'b00;
		14'h2b42: color = 2'b00;
		14'h2b43: color = 2'b00;
		14'h2b44: color = 2'b00;
		14'h2b45: color = 2'b00;
		14'h2b46: color = 2'b00;
		14'h2b47: color = 2'b00;
		14'h2b48: color = 2'b00;
		14'h2b49: color = 2'b00;
		14'h2b4a: color = 2'b00;
		14'h2b4b: color = 2'b00;
		14'h2b4c: color = 2'b00;
		14'h2b4d: color = 2'b00;
		14'h2b4e: color = 2'b00;
		14'h2b4f: color = 2'b00;
		14'h2b50: color = 2'b00;
		14'h2b51: color = 2'b00;
		14'h2b52: color = 2'b00;
		14'h2b53: color = 2'b00;
		14'h2b54: color = 2'b00;
		14'h2b55: color = 2'b00;
		14'h2b56: color = 2'b00;
		14'h2b57: color = 2'b00;
		14'h2b58: color = 2'b00;
		14'h2b59: color = 2'b00;
		14'h2b5a: color = 2'b01;
		14'h2b5b: color = 2'b11;
		14'h2b5c: color = 2'b11;
		14'h2b5d: color = 2'b11;
		14'h2b5e: color = 2'b11;
		14'h2b5f: color = 2'b11;
		14'h2b60: color = 2'b11;
		14'h2b61: color = 2'b11;
		14'h2b62: color = 2'b11;
		14'h2b63: color = 2'b11;
		14'h2b64: color = 2'b11;
		14'h2b65: color = 2'b11;
		14'h2b66: color = 2'b11;
		14'h2b67: color = 2'b11;
		14'h2b68: color = 2'b11;
		14'h2b69: color = 2'b11;
		14'h2b6a: color = 2'b11;
		14'h2b6b: color = 2'b11;
		14'h2b6c: color = 2'b11;
		14'h2b6d: color = 2'b11;
		14'h2b6e: color = 2'b11;
		14'h2b6f: color = 2'b11;
		14'h2b70: color = 2'b11;
		14'h2b71: color = 2'b11;
		14'h2b72: color = 2'b11;
		14'h2b73: color = 2'b11;
		14'h2b74: color = 2'b11;
		14'h2b75: color = 2'b11;
		14'h2b76: color = 2'b11;
		14'h2b77: color = 2'b11;
		14'h2b78: color = 2'b11;
		14'h2b79: color = 2'b11;
		14'h2b7a: color = 2'b11;
		14'h2b7b: color = 2'b11;
		14'h2b7c: color = 2'b11;
		14'h2b7d: color = 2'b11;
		14'h2b7e: color = 2'b11;
		14'h2b7f: color = 2'b11;
		14'h2b80: color = 2'b11;
		14'h2b81: color = 2'b11;
		14'h2b82: color = 2'b11;
		14'h2b83: color = 2'b11;
		14'h2b84: color = 2'b11;
		14'h2b85: color = 2'b11;
		14'h2b86: color = 2'b11;
		14'h2b87: color = 2'b11;
		14'h2b88: color = 2'b11;
		14'h2b89: color = 2'b11;
		14'h2b8a: color = 2'b11;
		14'h2b8b: color = 2'b11;
		14'h2b8c: color = 2'b11;
		14'h2b8d: color = 2'b11;
		14'h2b8e: color = 2'b11;
		14'h2b8f: color = 2'b11;
		14'h2b90: color = 2'b11;
		14'h2b91: color = 2'b11;
		14'h2b92: color = 2'b11;
		14'h2b93: color = 2'b11;
		14'h2b94: color = 2'b10;
		14'h2b95: color = 2'b01;
		14'h2b96: color = 2'b00;
		14'h2b97: color = 2'b00;
		14'h2b98: color = 2'b00;
		14'h2b99: color = 2'b00;
		14'h2b9a: color = 2'b01;
		14'h2b9b: color = 2'b00;
		14'h2b9c: color = 2'b00;
		14'h2b9d: color = 2'b00;
		14'h2b9e: color = 2'b00;
		14'h2b9f: color = 2'b00;
		14'h2ba0: color = 2'b00;
		14'h2ba1: color = 2'b00;
		14'h2ba2: color = 2'b01;
		14'h2ba3: color = 2'b00;
		14'h2ba4: color = 2'b01;
		14'h2ba5: color = 2'b00;
		14'h2ba6: color = 2'b00;
		14'h2ba7: color = 2'b00;
		14'h2ba8: color = 2'b00;
		14'h2ba9: color = 2'b00;
		14'h2baa: color = 2'b00;
		14'h2bab: color = 2'b00;
		14'h2bac: color = 2'b10;
		14'h2bad: color = 2'b11;
		14'h2bae: color = 2'b11;
		14'h2baf: color = 2'b11;
		14'h2bb0: color = 2'b11;
		14'h2bb1: color = 2'b11;
		14'h2bb2: color = 2'b10;
		14'h2bb3: color = 2'b10;
		14'h2bb4: color = 2'b10;
		14'h2bb5: color = 2'b01;
		14'h2bb6: color = 2'b00;
		14'h2bb7: color = 2'b00;
		14'h2bb8: color = 2'b00;
		14'h2bb9: color = 2'b00;
		14'h2bba: color = 2'b00;
		14'h2bbb: color = 2'b00;
		14'h2bbc: color = 2'b00;
		14'h2bbd: color = 2'b00;
		14'h2bbe: color = 2'b00;
		14'h2bbf: color = 2'b00;
		14'h2bc0: color = 2'b00;
		14'h2bc1: color = 2'b00;
		14'h2bc2: color = 2'b00;
		14'h2bc3: color = 2'b00;
		14'h2bc4: color = 2'b00;
		14'h2bc5: color = 2'b00;
		14'h2bc6: color = 2'b00;
		14'h2bc7: color = 2'b00;
		14'h2bc8: color = 2'b00;
		14'h2bc9: color = 2'b00;
		14'h2bca: color = 2'b00;
		14'h2bcb: color = 2'b00;
		14'h2bcc: color = 2'b00;
		14'h2bcd: color = 2'b00;
		14'h2bce: color = 2'b00;
		14'h2bcf: color = 2'b00;
		14'h2bd0: color = 2'b00;
		14'h2bd1: color = 2'b00;
		14'h2bd2: color = 2'b00;
		14'h2bd3: color = 2'b00;
		14'h2bd4: color = 2'b00;
		14'h2bd5: color = 2'b00;
		14'h2bd6: color = 2'b00;
		14'h2bd7: color = 2'b00;
		14'h2bd8: color = 2'b00;
		14'h2bd9: color = 2'b00;
		14'h2bda: color = 2'b00;
		14'h2bdb: color = 2'b01;
		14'h2bdc: color = 2'b01;
		14'h2bdd: color = 2'b10;
		14'h2bde: color = 2'b11;
		14'h2bdf: color = 2'b11;
		14'h2be0: color = 2'b11;
		14'h2be1: color = 2'b11;
		14'h2be2: color = 2'b11;
		14'h2be3: color = 2'b11;
		14'h2be4: color = 2'b11;
		14'h2be5: color = 2'b11;
		14'h2be6: color = 2'b11;
		14'h2be7: color = 2'b11;
		14'h2be8: color = 2'b11;
		14'h2be9: color = 2'b11;
		14'h2bea: color = 2'b11;
		14'h2beb: color = 2'b11;
		14'h2bec: color = 2'b11;
		14'h2bed: color = 2'b11;
		14'h2bee: color = 2'b11;
		14'h2bef: color = 2'b11;
		14'h2bf0: color = 2'b11;
		14'h2bf1: color = 2'b11;
		14'h2bf2: color = 2'b11;
		14'h2bf3: color = 2'b11;
		14'h2bf4: color = 2'b11;
		14'h2bf5: color = 2'b11;
		14'h2bf6: color = 2'b11;
		14'h2bf7: color = 2'b11;
		14'h2bf8: color = 2'b11;
		14'h2bf9: color = 2'b11;
		14'h2bfa: color = 2'b11;
		14'h2bfb: color = 2'b11;
		14'h2bfc: color = 2'b11;
		14'h2bfd: color = 2'b11;
		14'h2bfe: color = 2'b11;
		14'h2bff: color = 2'b11;
		14'h2c00: color = 2'b11;
		14'h2c01: color = 2'b11;
		14'h2c02: color = 2'b11;
		14'h2c03: color = 2'b11;
		14'h2c04: color = 2'b11;
		14'h2c05: color = 2'b11;
		14'h2c06: color = 2'b11;
		14'h2c07: color = 2'b11;
		14'h2c08: color = 2'b11;
		14'h2c09: color = 2'b11;
		14'h2c0a: color = 2'b11;
		14'h2c0b: color = 2'b11;
		14'h2c0c: color = 2'b11;
		14'h2c0d: color = 2'b11;
		14'h2c0e: color = 2'b11;
		14'h2c0f: color = 2'b11;
		14'h2c10: color = 2'b11;
		14'h2c11: color = 2'b11;
		14'h2c12: color = 2'b11;
		14'h2c13: color = 2'b11;
		14'h2c14: color = 2'b10;
		14'h2c15: color = 2'b01;
		14'h2c16: color = 2'b00;
		14'h2c17: color = 2'b00;
		14'h2c18: color = 2'b00;
		14'h2c19: color = 2'b00;
		14'h2c1a: color = 2'b01;
		14'h2c1b: color = 2'b00;
		14'h2c1c: color = 2'b00;
		14'h2c1d: color = 2'b00;
		14'h2c1e: color = 2'b00;
		14'h2c1f: color = 2'b00;
		14'h2c20: color = 2'b00;
		14'h2c21: color = 2'b00;
		14'h2c22: color = 2'b01;
		14'h2c23: color = 2'b00;
		14'h2c24: color = 2'b01;
		14'h2c25: color = 2'b00;
		14'h2c26: color = 2'b00;
		14'h2c27: color = 2'b00;
		14'h2c28: color = 2'b00;
		14'h2c29: color = 2'b00;
		14'h2c2a: color = 2'b00;
		14'h2c2b: color = 2'b00;
		14'h2c2c: color = 2'b10;
		14'h2c2d: color = 2'b11;
		14'h2c2e: color = 2'b11;
		14'h2c2f: color = 2'b11;
		14'h2c30: color = 2'b11;
		14'h2c31: color = 2'b11;
		14'h2c32: color = 2'b10;
		14'h2c33: color = 2'b10;
		14'h2c34: color = 2'b10;
		14'h2c35: color = 2'b01;
		14'h2c36: color = 2'b00;
		14'h2c37: color = 2'b00;
		14'h2c38: color = 2'b00;
		14'h2c39: color = 2'b00;
		14'h2c3a: color = 2'b00;
		14'h2c3b: color = 2'b00;
		14'h2c3c: color = 2'b00;
		14'h2c3d: color = 2'b00;
		14'h2c3e: color = 2'b00;
		14'h2c3f: color = 2'b00;
		14'h2c40: color = 2'b00;
		14'h2c41: color = 2'b00;
		14'h2c42: color = 2'b00;
		14'h2c43: color = 2'b00;
		14'h2c44: color = 2'b00;
		14'h2c45: color = 2'b00;
		14'h2c46: color = 2'b00;
		14'h2c47: color = 2'b00;
		14'h2c48: color = 2'b00;
		14'h2c49: color = 2'b00;
		14'h2c4a: color = 2'b00;
		14'h2c4b: color = 2'b00;
		14'h2c4c: color = 2'b00;
		14'h2c4d: color = 2'b00;
		14'h2c4e: color = 2'b00;
		14'h2c4f: color = 2'b00;
		14'h2c50: color = 2'b00;
		14'h2c51: color = 2'b00;
		14'h2c52: color = 2'b00;
		14'h2c53: color = 2'b00;
		14'h2c54: color = 2'b00;
		14'h2c55: color = 2'b00;
		14'h2c56: color = 2'b00;
		14'h2c57: color = 2'b00;
		14'h2c58: color = 2'b00;
		14'h2c59: color = 2'b00;
		14'h2c5a: color = 2'b00;
		14'h2c5b: color = 2'b01;
		14'h2c5c: color = 2'b01;
		14'h2c5d: color = 2'b10;
		14'h2c5e: color = 2'b11;
		14'h2c5f: color = 2'b11;
		14'h2c60: color = 2'b11;
		14'h2c61: color = 2'b11;
		14'h2c62: color = 2'b11;
		14'h2c63: color = 2'b11;
		14'h2c64: color = 2'b11;
		14'h2c65: color = 2'b11;
		14'h2c66: color = 2'b11;
		14'h2c67: color = 2'b11;
		14'h2c68: color = 2'b11;
		14'h2c69: color = 2'b11;
		14'h2c6a: color = 2'b11;
		14'h2c6b: color = 2'b11;
		14'h2c6c: color = 2'b11;
		14'h2c6d: color = 2'b11;
		14'h2c6e: color = 2'b11;
		14'h2c6f: color = 2'b11;
		14'h2c70: color = 2'b11;
		14'h2c71: color = 2'b11;
		14'h2c72: color = 2'b11;
		14'h2c73: color = 2'b11;
		14'h2c74: color = 2'b11;
		14'h2c75: color = 2'b11;
		14'h2c76: color = 2'b11;
		14'h2c77: color = 2'b11;
		14'h2c78: color = 2'b11;
		14'h2c79: color = 2'b11;
		14'h2c7a: color = 2'b11;
		14'h2c7b: color = 2'b11;
		14'h2c7c: color = 2'b11;
		14'h2c7d: color = 2'b11;
		14'h2c7e: color = 2'b11;
		14'h2c7f: color = 2'b11;
		14'h2c80: color = 2'b11;
		14'h2c81: color = 2'b11;
		14'h2c82: color = 2'b11;
		14'h2c83: color = 2'b11;
		14'h2c84: color = 2'b11;
		14'h2c85: color = 2'b11;
		14'h2c86: color = 2'b11;
		14'h2c87: color = 2'b11;
		14'h2c88: color = 2'b11;
		14'h2c89: color = 2'b11;
		14'h2c8a: color = 2'b11;
		14'h2c8b: color = 2'b11;
		14'h2c8c: color = 2'b11;
		14'h2c8d: color = 2'b11;
		14'h2c8e: color = 2'b11;
		14'h2c8f: color = 2'b11;
		14'h2c90: color = 2'b11;
		14'h2c91: color = 2'b11;
		14'h2c92: color = 2'b11;
		14'h2c93: color = 2'b01;
		14'h2c94: color = 2'b00;
		14'h2c95: color = 2'b00;
		14'h2c96: color = 2'b00;
		14'h2c97: color = 2'b00;
		14'h2c98: color = 2'b00;
		14'h2c99: color = 2'b00;
		14'h2c9a: color = 2'b00;
		14'h2c9b: color = 2'b00;
		14'h2c9c: color = 2'b00;
		14'h2c9d: color = 2'b00;
		14'h2c9e: color = 2'b00;
		14'h2c9f: color = 2'b00;
		14'h2ca0: color = 2'b00;
		14'h2ca1: color = 2'b00;
		14'h2ca2: color = 2'b00;
		14'h2ca3: color = 2'b00;
		14'h2ca4: color = 2'b01;
		14'h2ca5: color = 2'b01;
		14'h2ca6: color = 2'b00;
		14'h2ca7: color = 2'b01;
		14'h2ca8: color = 2'b01;
		14'h2ca9: color = 2'b00;
		14'h2caa: color = 2'b00;
		14'h2cab: color = 2'b00;
		14'h2cac: color = 2'b01;
		14'h2cad: color = 2'b11;
		14'h2cae: color = 2'b11;
		14'h2caf: color = 2'b11;
		14'h2cb0: color = 2'b11;
		14'h2cb1: color = 2'b11;
		14'h2cb2: color = 2'b10;
		14'h2cb3: color = 2'b10;
		14'h2cb4: color = 2'b10;
		14'h2cb5: color = 2'b10;
		14'h2cb6: color = 2'b01;
		14'h2cb7: color = 2'b01;
		14'h2cb8: color = 2'b01;
		14'h2cb9: color = 2'b00;
		14'h2cba: color = 2'b00;
		14'h2cbb: color = 2'b00;
		14'h2cbc: color = 2'b01;
		14'h2cbd: color = 2'b00;
		14'h2cbe: color = 2'b00;
		14'h2cbf: color = 2'b00;
		14'h2cc0: color = 2'b00;
		14'h2cc1: color = 2'b00;
		14'h2cc2: color = 2'b00;
		14'h2cc3: color = 2'b00;
		14'h2cc4: color = 2'b00;
		14'h2cc5: color = 2'b00;
		14'h2cc6: color = 2'b00;
		14'h2cc7: color = 2'b00;
		14'h2cc8: color = 2'b00;
		14'h2cc9: color = 2'b00;
		14'h2cca: color = 2'b00;
		14'h2ccb: color = 2'b00;
		14'h2ccc: color = 2'b00;
		14'h2ccd: color = 2'b00;
		14'h2cce: color = 2'b00;
		14'h2ccf: color = 2'b00;
		14'h2cd0: color = 2'b00;
		14'h2cd1: color = 2'b00;
		14'h2cd2: color = 2'b00;
		14'h2cd3: color = 2'b00;
		14'h2cd4: color = 2'b00;
		14'h2cd5: color = 2'b00;
		14'h2cd6: color = 2'b00;
		14'h2cd7: color = 2'b00;
		14'h2cd8: color = 2'b00;
		14'h2cd9: color = 2'b00;
		14'h2cda: color = 2'b00;
		14'h2cdb: color = 2'b00;
		14'h2cdc: color = 2'b00;
		14'h2cdd: color = 2'b00;
		14'h2cde: color = 2'b00;
		14'h2cdf: color = 2'b01;
		14'h2ce0: color = 2'b11;
		14'h2ce1: color = 2'b11;
		14'h2ce2: color = 2'b11;
		14'h2ce3: color = 2'b11;
		14'h2ce4: color = 2'b11;
		14'h2ce5: color = 2'b11;
		14'h2ce6: color = 2'b11;
		14'h2ce7: color = 2'b11;
		14'h2ce8: color = 2'b11;
		14'h2ce9: color = 2'b11;
		14'h2cea: color = 2'b11;
		14'h2ceb: color = 2'b11;
		14'h2cec: color = 2'b11;
		14'h2ced: color = 2'b11;
		14'h2cee: color = 2'b11;
		14'h2cef: color = 2'b11;
		14'h2cf0: color = 2'b11;
		14'h2cf1: color = 2'b11;
		14'h2cf2: color = 2'b11;
		14'h2cf3: color = 2'b11;
		14'h2cf4: color = 2'b11;
		14'h2cf5: color = 2'b11;
		14'h2cf6: color = 2'b11;
		14'h2cf7: color = 2'b11;
		14'h2cf8: color = 2'b11;
		14'h2cf9: color = 2'b11;
		14'h2cfa: color = 2'b11;
		14'h2cfb: color = 2'b11;
		14'h2cfc: color = 2'b11;
		14'h2cfd: color = 2'b11;
		14'h2cfe: color = 2'b11;
		14'h2cff: color = 2'b11;
		14'h2d00: color = 2'b11;
		14'h2d01: color = 2'b11;
		14'h2d02: color = 2'b11;
		14'h2d03: color = 2'b11;
		14'h2d04: color = 2'b11;
		14'h2d05: color = 2'b11;
		14'h2d06: color = 2'b11;
		14'h2d07: color = 2'b11;
		14'h2d08: color = 2'b11;
		14'h2d09: color = 2'b11;
		14'h2d0a: color = 2'b11;
		14'h2d0b: color = 2'b11;
		14'h2d0c: color = 2'b11;
		14'h2d0d: color = 2'b11;
		14'h2d0e: color = 2'b11;
		14'h2d0f: color = 2'b11;
		14'h2d10: color = 2'b11;
		14'h2d11: color = 2'b01;
		14'h2d12: color = 2'b01;
		14'h2d13: color = 2'b00;
		14'h2d14: color = 2'b00;
		14'h2d15: color = 2'b01;
		14'h2d16: color = 2'b00;
		14'h2d17: color = 2'b00;
		14'h2d18: color = 2'b00;
		14'h2d19: color = 2'b00;
		14'h2d1a: color = 2'b00;
		14'h2d1b: color = 2'b00;
		14'h2d1c: color = 2'b00;
		14'h2d1d: color = 2'b00;
		14'h2d1e: color = 2'b00;
		14'h2d1f: color = 2'b00;
		14'h2d20: color = 2'b00;
		14'h2d21: color = 2'b00;
		14'h2d22: color = 2'b00;
		14'h2d23: color = 2'b00;
		14'h2d24: color = 2'b01;
		14'h2d25: color = 2'b00;
		14'h2d26: color = 2'b00;
		14'h2d27: color = 2'b01;
		14'h2d28: color = 2'b01;
		14'h2d29: color = 2'b00;
		14'h2d2a: color = 2'b00;
		14'h2d2b: color = 2'b00;
		14'h2d2c: color = 2'b00;
		14'h2d2d: color = 2'b10;
		14'h2d2e: color = 2'b11;
		14'h2d2f: color = 2'b11;
		14'h2d30: color = 2'b11;
		14'h2d31: color = 2'b11;
		14'h2d32: color = 2'b11;
		14'h2d33: color = 2'b10;
		14'h2d34: color = 2'b10;
		14'h2d35: color = 2'b10;
		14'h2d36: color = 2'b10;
		14'h2d37: color = 2'b01;
		14'h2d38: color = 2'b01;
		14'h2d39: color = 2'b00;
		14'h2d3a: color = 2'b00;
		14'h2d3b: color = 2'b00;
		14'h2d3c: color = 2'b00;
		14'h2d3d: color = 2'b00;
		14'h2d3e: color = 2'b01;
		14'h2d3f: color = 2'b00;
		14'h2d40: color = 2'b00;
		14'h2d41: color = 2'b00;
		14'h2d42: color = 2'b00;
		14'h2d43: color = 2'b00;
		14'h2d44: color = 2'b00;
		14'h2d45: color = 2'b00;
		14'h2d46: color = 2'b00;
		14'h2d47: color = 2'b00;
		14'h2d48: color = 2'b00;
		14'h2d49: color = 2'b00;
		14'h2d4a: color = 2'b00;
		14'h2d4b: color = 2'b00;
		14'h2d4c: color = 2'b00;
		14'h2d4d: color = 2'b00;
		14'h2d4e: color = 2'b00;
		14'h2d4f: color = 2'b00;
		14'h2d50: color = 2'b00;
		14'h2d51: color = 2'b00;
		14'h2d52: color = 2'b00;
		14'h2d53: color = 2'b00;
		14'h2d54: color = 2'b00;
		14'h2d55: color = 2'b00;
		14'h2d56: color = 2'b00;
		14'h2d57: color = 2'b00;
		14'h2d58: color = 2'b00;
		14'h2d59: color = 2'b00;
		14'h2d5a: color = 2'b00;
		14'h2d5b: color = 2'b00;
		14'h2d5c: color = 2'b00;
		14'h2d5d: color = 2'b00;
		14'h2d5e: color = 2'b00;
		14'h2d5f: color = 2'b00;
		14'h2d60: color = 2'b00;
		14'h2d61: color = 2'b01;
		14'h2d62: color = 2'b11;
		14'h2d63: color = 2'b11;
		14'h2d64: color = 2'b11;
		14'h2d65: color = 2'b11;
		14'h2d66: color = 2'b11;
		14'h2d67: color = 2'b11;
		14'h2d68: color = 2'b11;
		14'h2d69: color = 2'b11;
		14'h2d6a: color = 2'b11;
		14'h2d6b: color = 2'b11;
		14'h2d6c: color = 2'b11;
		14'h2d6d: color = 2'b11;
		14'h2d6e: color = 2'b11;
		14'h2d6f: color = 2'b11;
		14'h2d70: color = 2'b11;
		14'h2d71: color = 2'b11;
		14'h2d72: color = 2'b11;
		14'h2d73: color = 2'b11;
		14'h2d74: color = 2'b11;
		14'h2d75: color = 2'b11;
		14'h2d76: color = 2'b11;
		14'h2d77: color = 2'b11;
		14'h2d78: color = 2'b11;
		14'h2d79: color = 2'b11;
		14'h2d7a: color = 2'b11;
		14'h2d7b: color = 2'b11;
		14'h2d7c: color = 2'b11;
		14'h2d7d: color = 2'b11;
		14'h2d7e: color = 2'b11;
		14'h2d7f: color = 2'b11;
		14'h2d80: color = 2'b11;
		14'h2d81: color = 2'b11;
		14'h2d82: color = 2'b11;
		14'h2d83: color = 2'b11;
		14'h2d84: color = 2'b11;
		14'h2d85: color = 2'b11;
		14'h2d86: color = 2'b11;
		14'h2d87: color = 2'b11;
		14'h2d88: color = 2'b11;
		14'h2d89: color = 2'b11;
		14'h2d8a: color = 2'b11;
		14'h2d8b: color = 2'b11;
		14'h2d8c: color = 2'b11;
		14'h2d8d: color = 2'b11;
		14'h2d8e: color = 2'b11;
		14'h2d8f: color = 2'b10;
		14'h2d90: color = 2'b00;
		14'h2d91: color = 2'b00;
		14'h2d92: color = 2'b01;
		14'h2d93: color = 2'b00;
		14'h2d94: color = 2'b00;
		14'h2d95: color = 2'b00;
		14'h2d96: color = 2'b00;
		14'h2d97: color = 2'b00;
		14'h2d98: color = 2'b00;
		14'h2d99: color = 2'b00;
		14'h2d9a: color = 2'b00;
		14'h2d9b: color = 2'b00;
		14'h2d9c: color = 2'b00;
		14'h2d9d: color = 2'b00;
		14'h2d9e: color = 2'b00;
		14'h2d9f: color = 2'b00;
		14'h2da0: color = 2'b00;
		14'h2da1: color = 2'b00;
		14'h2da2: color = 2'b00;
		14'h2da3: color = 2'b00;
		14'h2da4: color = 2'b00;
		14'h2da5: color = 2'b01;
		14'h2da6: color = 2'b00;
		14'h2da7: color = 2'b01;
		14'h2da8: color = 2'b01;
		14'h2da9: color = 2'b00;
		14'h2daa: color = 2'b01;
		14'h2dab: color = 2'b00;
		14'h2dac: color = 2'b00;
		14'h2dad: color = 2'b00;
		14'h2dae: color = 2'b11;
		14'h2daf: color = 2'b11;
		14'h2db0: color = 2'b11;
		14'h2db1: color = 2'b11;
		14'h2db2: color = 2'b11;
		14'h2db3: color = 2'b11;
		14'h2db4: color = 2'b10;
		14'h2db5: color = 2'b10;
		14'h2db6: color = 2'b10;
		14'h2db7: color = 2'b10;
		14'h2db8: color = 2'b10;
		14'h2db9: color = 2'b01;
		14'h2dba: color = 2'b00;
		14'h2dbb: color = 2'b00;
		14'h2dbc: color = 2'b00;
		14'h2dbd: color = 2'b00;
		14'h2dbe: color = 2'b00;
		14'h2dbf: color = 2'b00;
		14'h2dc0: color = 2'b00;
		14'h2dc1: color = 2'b00;
		14'h2dc2: color = 2'b00;
		14'h2dc3: color = 2'b00;
		14'h2dc4: color = 2'b00;
		14'h2dc5: color = 2'b00;
		14'h2dc6: color = 2'b00;
		14'h2dc7: color = 2'b00;
		14'h2dc8: color = 2'b00;
		14'h2dc9: color = 2'b00;
		14'h2dca: color = 2'b00;
		14'h2dcb: color = 2'b00;
		14'h2dcc: color = 2'b00;
		14'h2dcd: color = 2'b00;
		14'h2dce: color = 2'b00;
		14'h2dcf: color = 2'b00;
		14'h2dd0: color = 2'b00;
		14'h2dd1: color = 2'b00;
		14'h2dd2: color = 2'b00;
		14'h2dd3: color = 2'b00;
		14'h2dd4: color = 2'b00;
		14'h2dd5: color = 2'b00;
		14'h2dd6: color = 2'b00;
		14'h2dd7: color = 2'b00;
		14'h2dd8: color = 2'b00;
		14'h2dd9: color = 2'b00;
		14'h2dda: color = 2'b00;
		14'h2ddb: color = 2'b00;
		14'h2ddc: color = 2'b00;
		14'h2ddd: color = 2'b00;
		14'h2dde: color = 2'b00;
		14'h2ddf: color = 2'b00;
		14'h2de0: color = 2'b00;
		14'h2de1: color = 2'b00;
		14'h2de2: color = 2'b00;
		14'h2de3: color = 2'b01;
		14'h2de4: color = 2'b10;
		14'h2de5: color = 2'b11;
		14'h2de6: color = 2'b11;
		14'h2de7: color = 2'b11;
		14'h2de8: color = 2'b11;
		14'h2de9: color = 2'b11;
		14'h2dea: color = 2'b11;
		14'h2deb: color = 2'b11;
		14'h2dec: color = 2'b11;
		14'h2ded: color = 2'b11;
		14'h2dee: color = 2'b11;
		14'h2def: color = 2'b11;
		14'h2df0: color = 2'b11;
		14'h2df1: color = 2'b11;
		14'h2df2: color = 2'b11;
		14'h2df3: color = 2'b11;
		14'h2df4: color = 2'b11;
		14'h2df5: color = 2'b11;
		14'h2df6: color = 2'b11;
		14'h2df7: color = 2'b11;
		14'h2df8: color = 2'b11;
		14'h2df9: color = 2'b11;
		14'h2dfa: color = 2'b11;
		14'h2dfb: color = 2'b11;
		14'h2dfc: color = 2'b11;
		14'h2dfd: color = 2'b11;
		14'h2dfe: color = 2'b11;
		14'h2dff: color = 2'b11;
		14'h2e00: color = 2'b11;
		14'h2e01: color = 2'b11;
		14'h2e02: color = 2'b11;
		14'h2e03: color = 2'b11;
		14'h2e04: color = 2'b11;
		14'h2e05: color = 2'b11;
		14'h2e06: color = 2'b11;
		14'h2e07: color = 2'b11;
		14'h2e08: color = 2'b11;
		14'h2e09: color = 2'b11;
		14'h2e0a: color = 2'b11;
		14'h2e0b: color = 2'b11;
		14'h2e0c: color = 2'b11;
		14'h2e0d: color = 2'b10;
		14'h2e0e: color = 2'b01;
		14'h2e0f: color = 2'b01;
		14'h2e10: color = 2'b00;
		14'h2e11: color = 2'b01;
		14'h2e12: color = 2'b00;
		14'h2e13: color = 2'b00;
		14'h2e14: color = 2'b00;
		14'h2e15: color = 2'b01;
		14'h2e16: color = 2'b00;
		14'h2e17: color = 2'b00;
		14'h2e18: color = 2'b00;
		14'h2e19: color = 2'b00;
		14'h2e1a: color = 2'b00;
		14'h2e1b: color = 2'b00;
		14'h2e1c: color = 2'b00;
		14'h2e1d: color = 2'b00;
		14'h2e1e: color = 2'b00;
		14'h2e1f: color = 2'b00;
		14'h2e20: color = 2'b00;
		14'h2e21: color = 2'b00;
		14'h2e22: color = 2'b00;
		14'h2e23: color = 2'b00;
		14'h2e24: color = 2'b00;
		14'h2e25: color = 2'b01;
		14'h2e26: color = 2'b00;
		14'h2e27: color = 2'b01;
		14'h2e28: color = 2'b01;
		14'h2e29: color = 2'b00;
		14'h2e2a: color = 2'b00;
		14'h2e2b: color = 2'b00;
		14'h2e2c: color = 2'b00;
		14'h2e2d: color = 2'b00;
		14'h2e2e: color = 2'b10;
		14'h2e2f: color = 2'b11;
		14'h2e30: color = 2'b11;
		14'h2e31: color = 2'b11;
		14'h2e32: color = 2'b11;
		14'h2e33: color = 2'b11;
		14'h2e34: color = 2'b10;
		14'h2e35: color = 2'b10;
		14'h2e36: color = 2'b10;
		14'h2e37: color = 2'b10;
		14'h2e38: color = 2'b10;
		14'h2e39: color = 2'b10;
		14'h2e3a: color = 2'b01;
		14'h2e3b: color = 2'b00;
		14'h2e3c: color = 2'b00;
		14'h2e3d: color = 2'b00;
		14'h2e3e: color = 2'b00;
		14'h2e3f: color = 2'b00;
		14'h2e40: color = 2'b00;
		14'h2e41: color = 2'b00;
		14'h2e42: color = 2'b00;
		14'h2e43: color = 2'b00;
		14'h2e44: color = 2'b00;
		14'h2e45: color = 2'b00;
		14'h2e46: color = 2'b00;
		14'h2e47: color = 2'b00;
		14'h2e48: color = 2'b00;
		14'h2e49: color = 2'b00;
		14'h2e4a: color = 2'b00;
		14'h2e4b: color = 2'b00;
		14'h2e4c: color = 2'b00;
		14'h2e4d: color = 2'b00;
		14'h2e4e: color = 2'b00;
		14'h2e4f: color = 2'b00;
		14'h2e50: color = 2'b00;
		14'h2e51: color = 2'b00;
		14'h2e52: color = 2'b00;
		14'h2e53: color = 2'b00;
		14'h2e54: color = 2'b00;
		14'h2e55: color = 2'b00;
		14'h2e56: color = 2'b00;
		14'h2e57: color = 2'b00;
		14'h2e58: color = 2'b00;
		14'h2e59: color = 2'b00;
		14'h2e5a: color = 2'b00;
		14'h2e5b: color = 2'b00;
		14'h2e5c: color = 2'b00;
		14'h2e5d: color = 2'b00;
		14'h2e5e: color = 2'b00;
		14'h2e5f: color = 2'b00;
		14'h2e60: color = 2'b00;
		14'h2e61: color = 2'b00;
		14'h2e62: color = 2'b00;
		14'h2e63: color = 2'b00;
		14'h2e64: color = 2'b00;
		14'h2e65: color = 2'b00;
		14'h2e66: color = 2'b01;
		14'h2e67: color = 2'b11;
		14'h2e68: color = 2'b11;
		14'h2e69: color = 2'b11;
		14'h2e6a: color = 2'b11;
		14'h2e6b: color = 2'b11;
		14'h2e6c: color = 2'b11;
		14'h2e6d: color = 2'b11;
		14'h2e6e: color = 2'b11;
		14'h2e6f: color = 2'b11;
		14'h2e70: color = 2'b11;
		14'h2e71: color = 2'b11;
		14'h2e72: color = 2'b11;
		14'h2e73: color = 2'b11;
		14'h2e74: color = 2'b11;
		14'h2e75: color = 2'b11;
		14'h2e76: color = 2'b11;
		14'h2e77: color = 2'b11;
		14'h2e78: color = 2'b11;
		14'h2e79: color = 2'b11;
		14'h2e7a: color = 2'b11;
		14'h2e7b: color = 2'b11;
		14'h2e7c: color = 2'b11;
		14'h2e7d: color = 2'b11;
		14'h2e7e: color = 2'b11;
		14'h2e7f: color = 2'b11;
		14'h2e80: color = 2'b11;
		14'h2e81: color = 2'b11;
		14'h2e82: color = 2'b11;
		14'h2e83: color = 2'b11;
		14'h2e84: color = 2'b11;
		14'h2e85: color = 2'b11;
		14'h2e86: color = 2'b11;
		14'h2e87: color = 2'b11;
		14'h2e88: color = 2'b11;
		14'h2e89: color = 2'b11;
		14'h2e8a: color = 2'b11;
		14'h2e8b: color = 2'b10;
		14'h2e8c: color = 2'b01;
		14'h2e8d: color = 2'b00;
		14'h2e8e: color = 2'b00;
		14'h2e8f: color = 2'b00;
		14'h2e90: color = 2'b00;
		14'h2e91: color = 2'b00;
		14'h2e92: color = 2'b00;
		14'h2e93: color = 2'b01;
		14'h2e94: color = 2'b00;
		14'h2e95: color = 2'b00;
		14'h2e96: color = 2'b00;
		14'h2e97: color = 2'b01;
		14'h2e98: color = 2'b01;
		14'h2e99: color = 2'b00;
		14'h2e9a: color = 2'b00;
		14'h2e9b: color = 2'b00;
		14'h2e9c: color = 2'b00;
		14'h2e9d: color = 2'b00;
		14'h2e9e: color = 2'b00;
		14'h2e9f: color = 2'b00;
		14'h2ea0: color = 2'b00;
		14'h2ea1: color = 2'b00;
		14'h2ea2: color = 2'b00;
		14'h2ea3: color = 2'b00;
		14'h2ea4: color = 2'b00;
		14'h2ea5: color = 2'b00;
		14'h2ea6: color = 2'b01;
		14'h2ea7: color = 2'b00;
		14'h2ea8: color = 2'b00;
		14'h2ea9: color = 2'b00;
		14'h2eaa: color = 2'b00;
		14'h2eab: color = 2'b00;
		14'h2eac: color = 2'b00;
		14'h2ead: color = 2'b00;
		14'h2eae: color = 2'b00;
		14'h2eaf: color = 2'b11;
		14'h2eb0: color = 2'b11;
		14'h2eb1: color = 2'b11;
		14'h2eb2: color = 2'b11;
		14'h2eb3: color = 2'b11;
		14'h2eb4: color = 2'b11;
		14'h2eb5: color = 2'b10;
		14'h2eb6: color = 2'b10;
		14'h2eb7: color = 2'b10;
		14'h2eb8: color = 2'b10;
		14'h2eb9: color = 2'b01;
		14'h2eba: color = 2'b01;
		14'h2ebb: color = 2'b01;
		14'h2ebc: color = 2'b01;
		14'h2ebd: color = 2'b00;
		14'h2ebe: color = 2'b00;
		14'h2ebf: color = 2'b00;
		14'h2ec0: color = 2'b00;
		14'h2ec1: color = 2'b00;
		14'h2ec2: color = 2'b00;
		14'h2ec3: color = 2'b00;
		14'h2ec4: color = 2'b00;
		14'h2ec5: color = 2'b00;
		14'h2ec6: color = 2'b00;
		14'h2ec7: color = 2'b00;
		14'h2ec8: color = 2'b00;
		14'h2ec9: color = 2'b00;
		14'h2eca: color = 2'b00;
		14'h2ecb: color = 2'b00;
		14'h2ecc: color = 2'b00;
		14'h2ecd: color = 2'b00;
		14'h2ece: color = 2'b00;
		14'h2ecf: color = 2'b00;
		14'h2ed0: color = 2'b00;
		14'h2ed1: color = 2'b00;
		14'h2ed2: color = 2'b00;
		14'h2ed3: color = 2'b00;
		14'h2ed4: color = 2'b00;
		14'h2ed5: color = 2'b00;
		14'h2ed6: color = 2'b00;
		14'h2ed7: color = 2'b00;
		14'h2ed8: color = 2'b00;
		14'h2ed9: color = 2'b00;
		14'h2eda: color = 2'b00;
		14'h2edb: color = 2'b00;
		14'h2edc: color = 2'b00;
		14'h2edd: color = 2'b00;
		14'h2ede: color = 2'b00;
		14'h2edf: color = 2'b00;
		14'h2ee0: color = 2'b00;
		14'h2ee1: color = 2'b00;
		14'h2ee2: color = 2'b00;
		14'h2ee3: color = 2'b00;
		14'h2ee4: color = 2'b00;
		14'h2ee5: color = 2'b00;
		14'h2ee6: color = 2'b00;
		14'h2ee7: color = 2'b00;
		14'h2ee8: color = 2'b00;
		14'h2ee9: color = 2'b10;
		14'h2eea: color = 2'b11;
		14'h2eeb: color = 2'b11;
		14'h2eec: color = 2'b11;
		14'h2eed: color = 2'b11;
		14'h2eee: color = 2'b11;
		14'h2eef: color = 2'b11;
		14'h2ef0: color = 2'b11;
		14'h2ef1: color = 2'b11;
		14'h2ef2: color = 2'b11;
		14'h2ef3: color = 2'b11;
		14'h2ef4: color = 2'b11;
		14'h2ef5: color = 2'b11;
		14'h2ef6: color = 2'b11;
		14'h2ef7: color = 2'b11;
		14'h2ef8: color = 2'b11;
		14'h2ef9: color = 2'b11;
		14'h2efa: color = 2'b11;
		14'h2efb: color = 2'b11;
		14'h2efc: color = 2'b11;
		14'h2efd: color = 2'b11;
		14'h2efe: color = 2'b11;
		14'h2eff: color = 2'b11;
		14'h2f00: color = 2'b11;
		14'h2f01: color = 2'b11;
		14'h2f02: color = 2'b11;
		14'h2f03: color = 2'b11;
		14'h2f04: color = 2'b11;
		14'h2f05: color = 2'b11;
		14'h2f06: color = 2'b11;
		14'h2f07: color = 2'b11;
		14'h2f08: color = 2'b11;
		14'h2f09: color = 2'b01;
		14'h2f0a: color = 2'b01;
		14'h2f0b: color = 2'b00;
		14'h2f0c: color = 2'b00;
		14'h2f0d: color = 2'b01;
		14'h2f0e: color = 2'b01;
		14'h2f0f: color = 2'b00;
		14'h2f10: color = 2'b01;
		14'h2f11: color = 2'b00;
		14'h2f12: color = 2'b00;
		14'h2f13: color = 2'b00;
		14'h2f14: color = 2'b00;
		14'h2f15: color = 2'b00;
		14'h2f16: color = 2'b00;
		14'h2f17: color = 2'b00;
		14'h2f18: color = 2'b00;
		14'h2f19: color = 2'b00;
		14'h2f1a: color = 2'b00;
		14'h2f1b: color = 2'b00;
		14'h2f1c: color = 2'b00;
		14'h2f1d: color = 2'b00;
		14'h2f1e: color = 2'b00;
		14'h2f1f: color = 2'b00;
		14'h2f20: color = 2'b00;
		14'h2f21: color = 2'b00;
		14'h2f22: color = 2'b00;
		14'h2f23: color = 2'b01;
		14'h2f24: color = 2'b00;
		14'h2f25: color = 2'b01;
		14'h2f26: color = 2'b01;
		14'h2f27: color = 2'b00;
		14'h2f28: color = 2'b00;
		14'h2f29: color = 2'b01;
		14'h2f2a: color = 2'b00;
		14'h2f2b: color = 2'b00;
		14'h2f2c: color = 2'b00;
		14'h2f2d: color = 2'b00;
		14'h2f2e: color = 2'b00;
		14'h2f2f: color = 2'b01;
		14'h2f30: color = 2'b11;
		14'h2f31: color = 2'b11;
		14'h2f32: color = 2'b11;
		14'h2f33: color = 2'b11;
		14'h2f34: color = 2'b11;
		14'h2f35: color = 2'b11;
		14'h2f36: color = 2'b10;
		14'h2f37: color = 2'b10;
		14'h2f38: color = 2'b10;
		14'h2f39: color = 2'b10;
		14'h2f3a: color = 2'b10;
		14'h2f3b: color = 2'b10;
		14'h2f3c: color = 2'b01;
		14'h2f3d: color = 2'b01;
		14'h2f3e: color = 2'b01;
		14'h2f3f: color = 2'b00;
		14'h2f40: color = 2'b01;
		14'h2f41: color = 2'b00;
		14'h2f42: color = 2'b00;
		14'h2f43: color = 2'b00;
		14'h2f44: color = 2'b00;
		14'h2f45: color = 2'b00;
		14'h2f46: color = 2'b00;
		14'h2f47: color = 2'b00;
		14'h2f48: color = 2'b00;
		14'h2f49: color = 2'b00;
		14'h2f4a: color = 2'b00;
		14'h2f4b: color = 2'b00;
		14'h2f4c: color = 2'b00;
		14'h2f4d: color = 2'b00;
		14'h2f4e: color = 2'b00;
		14'h2f4f: color = 2'b00;
		14'h2f50: color = 2'b00;
		14'h2f51: color = 2'b00;
		14'h2f52: color = 2'b00;
		14'h2f53: color = 2'b00;
		14'h2f54: color = 2'b00;
		14'h2f55: color = 2'b00;
		14'h2f56: color = 2'b00;
		14'h2f57: color = 2'b00;
		14'h2f58: color = 2'b00;
		14'h2f59: color = 2'b00;
		14'h2f5a: color = 2'b00;
		14'h2f5b: color = 2'b00;
		14'h2f5c: color = 2'b00;
		14'h2f5d: color = 2'b00;
		14'h2f5e: color = 2'b00;
		14'h2f5f: color = 2'b00;
		14'h2f60: color = 2'b00;
		14'h2f61: color = 2'b00;
		14'h2f62: color = 2'b00;
		14'h2f63: color = 2'b00;
		14'h2f64: color = 2'b00;
		14'h2f65: color = 2'b00;
		14'h2f66: color = 2'b00;
		14'h2f67: color = 2'b00;
		14'h2f68: color = 2'b00;
		14'h2f69: color = 2'b00;
		14'h2f6a: color = 2'b00;
		14'h2f6b: color = 2'b10;
		14'h2f6c: color = 2'b11;
		14'h2f6d: color = 2'b11;
		14'h2f6e: color = 2'b11;
		14'h2f6f: color = 2'b11;
		14'h2f70: color = 2'b11;
		14'h2f71: color = 2'b11;
		14'h2f72: color = 2'b11;
		14'h2f73: color = 2'b11;
		14'h2f74: color = 2'b11;
		14'h2f75: color = 2'b11;
		14'h2f76: color = 2'b11;
		14'h2f77: color = 2'b11;
		14'h2f78: color = 2'b11;
		14'h2f79: color = 2'b11;
		14'h2f7a: color = 2'b11;
		14'h2f7b: color = 2'b11;
		14'h2f7c: color = 2'b11;
		14'h2f7d: color = 2'b11;
		14'h2f7e: color = 2'b11;
		14'h2f7f: color = 2'b11;
		14'h2f80: color = 2'b11;
		14'h2f81: color = 2'b11;
		14'h2f82: color = 2'b11;
		14'h2f83: color = 2'b11;
		14'h2f84: color = 2'b11;
		14'h2f85: color = 2'b11;
		14'h2f86: color = 2'b10;
		14'h2f87: color = 2'b01;
		14'h2f88: color = 2'b01;
		14'h2f89: color = 2'b00;
		14'h2f8a: color = 2'b01;
		14'h2f8b: color = 2'b00;
		14'h2f8c: color = 2'b01;
		14'h2f8d: color = 2'b00;
		14'h2f8e: color = 2'b00;
		14'h2f8f: color = 2'b00;
		14'h2f90: color = 2'b00;
		14'h2f91: color = 2'b00;
		14'h2f92: color = 2'b01;
		14'h2f93: color = 2'b00;
		14'h2f94: color = 2'b00;
		14'h2f95: color = 2'b00;
		14'h2f96: color = 2'b00;
		14'h2f97: color = 2'b00;
		14'h2f98: color = 2'b00;
		14'h2f99: color = 2'b00;
		14'h2f9a: color = 2'b00;
		14'h2f9b: color = 2'b00;
		14'h2f9c: color = 2'b00;
		14'h2f9d: color = 2'b00;
		14'h2f9e: color = 2'b00;
		14'h2f9f: color = 2'b00;
		14'h2fa0: color = 2'b00;
		14'h2fa1: color = 2'b00;
		14'h2fa2: color = 2'b00;
		14'h2fa3: color = 2'b00;
		14'h2fa4: color = 2'b00;
		14'h2fa5: color = 2'b00;
		14'h2fa6: color = 2'b00;
		14'h2fa7: color = 2'b00;
		14'h2fa8: color = 2'b00;
		14'h2fa9: color = 2'b01;
		14'h2faa: color = 2'b00;
		14'h2fab: color = 2'b01;
		14'h2fac: color = 2'b00;
		14'h2fad: color = 2'b00;
		14'h2fae: color = 2'b00;
		14'h2faf: color = 2'b01;
		14'h2fb0: color = 2'b11;
		14'h2fb1: color = 2'b11;
		14'h2fb2: color = 2'b11;
		14'h2fb3: color = 2'b11;
		14'h2fb4: color = 2'b11;
		14'h2fb5: color = 2'b11;
		14'h2fb6: color = 2'b11;
		14'h2fb7: color = 2'b10;
		14'h2fb8: color = 2'b10;
		14'h2fb9: color = 2'b01;
		14'h2fba: color = 2'b10;
		14'h2fbb: color = 2'b01;
		14'h2fbc: color = 2'b10;
		14'h2fbd: color = 2'b01;
		14'h2fbe: color = 2'b01;
		14'h2fbf: color = 2'b00;
		14'h2fc0: color = 2'b00;
		14'h2fc1: color = 2'b00;
		14'h2fc2: color = 2'b00;
		14'h2fc3: color = 2'b00;
		14'h2fc4: color = 2'b00;
		14'h2fc5: color = 2'b00;
		14'h2fc6: color = 2'b00;
		14'h2fc7: color = 2'b00;
		14'h2fc8: color = 2'b00;
		14'h2fc9: color = 2'b00;
		14'h2fca: color = 2'b00;
		14'h2fcb: color = 2'b00;
		14'h2fcc: color = 2'b00;
		14'h2fcd: color = 2'b00;
		14'h2fce: color = 2'b00;
		14'h2fcf: color = 2'b00;
		14'h2fd0: color = 2'b00;
		14'h2fd1: color = 2'b00;
		14'h2fd2: color = 2'b00;
		14'h2fd3: color = 2'b00;
		14'h2fd4: color = 2'b00;
		14'h2fd5: color = 2'b00;
		14'h2fd6: color = 2'b00;
		14'h2fd7: color = 2'b00;
		14'h2fd8: color = 2'b00;
		14'h2fd9: color = 2'b00;
		14'h2fda: color = 2'b00;
		14'h2fdb: color = 2'b00;
		14'h2fdc: color = 2'b00;
		14'h2fdd: color = 2'b00;
		14'h2fde: color = 2'b00;
		14'h2fdf: color = 2'b00;
		14'h2fe0: color = 2'b00;
		14'h2fe1: color = 2'b00;
		14'h2fe2: color = 2'b00;
		14'h2fe3: color = 2'b00;
		14'h2fe4: color = 2'b00;
		14'h2fe5: color = 2'b00;
		14'h2fe6: color = 2'b00;
		14'h2fe7: color = 2'b00;
		14'h2fe8: color = 2'b00;
		14'h2fe9: color = 2'b00;
		14'h2fea: color = 2'b00;
		14'h2feb: color = 2'b00;
		14'h2fec: color = 2'b00;
		14'h2fed: color = 2'b11;
		14'h2fee: color = 2'b11;
		14'h2fef: color = 2'b11;
		14'h2ff0: color = 2'b11;
		14'h2ff1: color = 2'b11;
		14'h2ff2: color = 2'b11;
		14'h2ff3: color = 2'b11;
		14'h2ff4: color = 2'b11;
		14'h2ff5: color = 2'b11;
		14'h2ff6: color = 2'b11;
		14'h2ff7: color = 2'b11;
		14'h2ff8: color = 2'b11;
		14'h2ff9: color = 2'b11;
		14'h2ffa: color = 2'b11;
		14'h2ffb: color = 2'b11;
		14'h2ffc: color = 2'b11;
		14'h2ffd: color = 2'b11;
		14'h2ffe: color = 2'b11;
		14'h2fff: color = 2'b11;
		14'h3000: color = 2'b11;
		14'h3001: color = 2'b11;
		14'h3002: color = 2'b11;
		14'h3003: color = 2'b10;
		14'h3004: color = 2'b01;
		14'h3005: color = 2'b10;
		14'h3006: color = 2'b01;
		14'h3007: color = 2'b00;
		14'h3008: color = 2'b00;
		14'h3009: color = 2'b00;
		14'h300a: color = 2'b01;
		14'h300b: color = 2'b00;
		14'h300c: color = 2'b00;
		14'h300d: color = 2'b00;
		14'h300e: color = 2'b01;
		14'h300f: color = 2'b00;
		14'h3010: color = 2'b01;
		14'h3011: color = 2'b00;
		14'h3012: color = 2'b00;
		14'h3013: color = 2'b00;
		14'h3014: color = 2'b00;
		14'h3015: color = 2'b00;
		14'h3016: color = 2'b00;
		14'h3017: color = 2'b00;
		14'h3018: color = 2'b00;
		14'h3019: color = 2'b00;
		14'h301a: color = 2'b00;
		14'h301b: color = 2'b00;
		14'h301c: color = 2'b00;
		14'h301d: color = 2'b00;
		14'h301e: color = 2'b00;
		14'h301f: color = 2'b00;
		14'h3020: color = 2'b00;
		14'h3021: color = 2'b00;
		14'h3022: color = 2'b00;
		14'h3023: color = 2'b00;
		14'h3024: color = 2'b00;
		14'h3025: color = 2'b00;
		14'h3026: color = 2'b01;
		14'h3027: color = 2'b00;
		14'h3028: color = 2'b00;
		14'h3029: color = 2'b01;
		14'h302a: color = 2'b00;
		14'h302b: color = 2'b00;
		14'h302c: color = 2'b00;
		14'h302d: color = 2'b00;
		14'h302e: color = 2'b00;
		14'h302f: color = 2'b00;
		14'h3030: color = 2'b01;
		14'h3031: color = 2'b11;
		14'h3032: color = 2'b11;
		14'h3033: color = 2'b11;
		14'h3034: color = 2'b11;
		14'h3035: color = 2'b11;
		14'h3036: color = 2'b11;
		14'h3037: color = 2'b11;
		14'h3038: color = 2'b11;
		14'h3039: color = 2'b10;
		14'h303a: color = 2'b10;
		14'h303b: color = 2'b10;
		14'h303c: color = 2'b01;
		14'h303d: color = 2'b10;
		14'h303e: color = 2'b01;
		14'h303f: color = 2'b01;
		14'h3040: color = 2'b01;
		14'h3041: color = 2'b01;
		14'h3042: color = 2'b00;
		14'h3043: color = 2'b00;
		14'h3044: color = 2'b00;
		14'h3045: color = 2'b00;
		14'h3046: color = 2'b00;
		14'h3047: color = 2'b00;
		14'h3048: color = 2'b00;
		14'h3049: color = 2'b00;
		14'h304a: color = 2'b00;
		14'h304b: color = 2'b00;
		14'h304c: color = 2'b00;
		14'h304d: color = 2'b00;
		14'h304e: color = 2'b00;
		14'h304f: color = 2'b00;
		14'h3050: color = 2'b00;
		14'h3051: color = 2'b00;
		14'h3052: color = 2'b00;
		14'h3053: color = 2'b00;
		14'h3054: color = 2'b00;
		14'h3055: color = 2'b00;
		14'h3056: color = 2'b00;
		14'h3057: color = 2'b00;
		14'h3058: color = 2'b00;
		14'h3059: color = 2'b00;
		14'h305a: color = 2'b00;
		14'h305b: color = 2'b00;
		14'h305c: color = 2'b00;
		14'h305d: color = 2'b00;
		14'h305e: color = 2'b00;
		14'h305f: color = 2'b00;
		14'h3060: color = 2'b00;
		14'h3061: color = 2'b00;
		14'h3062: color = 2'b00;
		14'h3063: color = 2'b00;
		14'h3064: color = 2'b00;
		14'h3065: color = 2'b00;
		14'h3066: color = 2'b00;
		14'h3067: color = 2'b00;
		14'h3068: color = 2'b00;
		14'h3069: color = 2'b00;
		14'h306a: color = 2'b00;
		14'h306b: color = 2'b00;
		14'h306c: color = 2'b00;
		14'h306d: color = 2'b00;
		14'h306e: color = 2'b01;
		14'h306f: color = 2'b11;
		14'h3070: color = 2'b11;
		14'h3071: color = 2'b11;
		14'h3072: color = 2'b11;
		14'h3073: color = 2'b11;
		14'h3074: color = 2'b11;
		14'h3075: color = 2'b11;
		14'h3076: color = 2'b11;
		14'h3077: color = 2'b11;
		14'h3078: color = 2'b11;
		14'h3079: color = 2'b11;
		14'h307a: color = 2'b11;
		14'h307b: color = 2'b11;
		14'h307c: color = 2'b11;
		14'h307d: color = 2'b11;
		14'h307e: color = 2'b11;
		14'h307f: color = 2'b11;
		14'h3080: color = 2'b11;
		14'h3081: color = 2'b10;
		14'h3082: color = 2'b10;
		14'h3083: color = 2'b01;
		14'h3084: color = 2'b01;
		14'h3085: color = 2'b00;
		14'h3086: color = 2'b01;
		14'h3087: color = 2'b00;
		14'h3088: color = 2'b00;
		14'h3089: color = 2'b00;
		14'h308a: color = 2'b01;
		14'h308b: color = 2'b00;
		14'h308c: color = 2'b01;
		14'h308d: color = 2'b00;
		14'h308e: color = 2'b00;
		14'h308f: color = 2'b00;
		14'h3090: color = 2'b00;
		14'h3091: color = 2'b00;
		14'h3092: color = 2'b00;
		14'h3093: color = 2'b01;
		14'h3094: color = 2'b00;
		14'h3095: color = 2'b00;
		14'h3096: color = 2'b00;
		14'h3097: color = 2'b00;
		14'h3098: color = 2'b00;
		14'h3099: color = 2'b00;
		14'h309a: color = 2'b00;
		14'h309b: color = 2'b00;
		14'h309c: color = 2'b00;
		14'h309d: color = 2'b00;
		14'h309e: color = 2'b00;
		14'h309f: color = 2'b00;
		14'h30a0: color = 2'b00;
		14'h30a1: color = 2'b00;
		14'h30a2: color = 2'b00;
		14'h30a3: color = 2'b00;
		14'h30a4: color = 2'b00;
		14'h30a5: color = 2'b00;
		14'h30a6: color = 2'b00;
		14'h30a7: color = 2'b00;
		14'h30a8: color = 2'b00;
		14'h30a9: color = 2'b00;
		14'h30aa: color = 2'b00;
		14'h30ab: color = 2'b00;
		14'h30ac: color = 2'b00;
		14'h30ad: color = 2'b00;
		14'h30ae: color = 2'b00;
		14'h30af: color = 2'b00;
		14'h30b0: color = 2'b00;
		14'h30b1: color = 2'b11;
		14'h30b2: color = 2'b11;
		14'h30b3: color = 2'b11;
		14'h30b4: color = 2'b11;
		14'h30b5: color = 2'b11;
		14'h30b6: color = 2'b11;
		14'h30b7: color = 2'b11;
		14'h30b8: color = 2'b11;
		14'h30b9: color = 2'b11;
		14'h30ba: color = 2'b10;
		14'h30bb: color = 2'b01;
		14'h30bc: color = 2'b01;
		14'h30bd: color = 2'b01;
		14'h30be: color = 2'b01;
		14'h30bf: color = 2'b01;
		14'h30c0: color = 2'b01;
		14'h30c1: color = 2'b01;
		14'h30c2: color = 2'b01;
		14'h30c3: color = 2'b00;
		14'h30c4: color = 2'b00;
		14'h30c5: color = 2'b00;
		14'h30c6: color = 2'b00;
		14'h30c7: color = 2'b00;
		14'h30c8: color = 2'b00;
		14'h30c9: color = 2'b00;
		14'h30ca: color = 2'b00;
		14'h30cb: color = 2'b00;
		14'h30cc: color = 2'b00;
		14'h30cd: color = 2'b00;
		14'h30ce: color = 2'b00;
		14'h30cf: color = 2'b00;
		14'h30d0: color = 2'b10;
		14'h30d1: color = 2'b01;
		14'h30d2: color = 2'b00;
		14'h30d3: color = 2'b00;
		14'h30d4: color = 2'b00;
		14'h30d5: color = 2'b00;
		14'h30d6: color = 2'b00;
		14'h30d7: color = 2'b00;
		14'h30d8: color = 2'b00;
		14'h30d9: color = 2'b00;
		14'h30da: color = 2'b00;
		14'h30db: color = 2'b00;
		14'h30dc: color = 2'b00;
		14'h30dd: color = 2'b00;
		14'h30de: color = 2'b00;
		14'h30df: color = 2'b00;
		14'h30e0: color = 2'b00;
		14'h30e1: color = 2'b00;
		14'h30e2: color = 2'b00;
		14'h30e3: color = 2'b00;
		14'h30e4: color = 2'b00;
		14'h30e5: color = 2'b00;
		14'h30e6: color = 2'b00;
		14'h30e7: color = 2'b00;
		14'h30e8: color = 2'b00;
		14'h30e9: color = 2'b00;
		14'h30ea: color = 2'b00;
		14'h30eb: color = 2'b00;
		14'h30ec: color = 2'b00;
		14'h30ed: color = 2'b00;
		14'h30ee: color = 2'b00;
		14'h30ef: color = 2'b00;
		14'h30f0: color = 2'b11;
		14'h30f1: color = 2'b11;
		14'h30f2: color = 2'b11;
		14'h30f3: color = 2'b11;
		14'h30f4: color = 2'b11;
		14'h30f5: color = 2'b11;
		14'h30f6: color = 2'b11;
		14'h30f7: color = 2'b11;
		14'h30f8: color = 2'b11;
		14'h30f9: color = 2'b11;
		14'h30fa: color = 2'b11;
		14'h30fb: color = 2'b11;
		14'h30fc: color = 2'b11;
		14'h30fd: color = 2'b11;
		14'h30fe: color = 2'b11;
		14'h30ff: color = 2'b11;
		14'h3100: color = 2'b00;
		14'h3101: color = 2'b10;
		14'h3102: color = 2'b00;
		14'h3103: color = 2'b01;
		14'h3104: color = 2'b00;
		14'h3105: color = 2'b00;
		14'h3106: color = 2'b00;
		14'h3107: color = 2'b01;
		14'h3108: color = 2'b01;
		14'h3109: color = 2'b00;
		14'h310a: color = 2'b01;
		14'h310b: color = 2'b00;
		14'h310c: color = 2'b00;
		14'h310d: color = 2'b01;
		14'h310e: color = 2'b00;
		14'h310f: color = 2'b00;
		14'h3110: color = 2'b00;
		14'h3111: color = 2'b01;
		14'h3112: color = 2'b00;
		14'h3113: color = 2'b00;
		14'h3114: color = 2'b00;
		14'h3115: color = 2'b00;
		14'h3116: color = 2'b00;
		14'h3117: color = 2'b00;
		14'h3118: color = 2'b00;
		14'h3119: color = 2'b00;
		14'h311a: color = 2'b00;
		14'h311b: color = 2'b00;
		14'h311c: color = 2'b00;
		14'h311d: color = 2'b00;
		14'h311e: color = 2'b00;
		14'h311f: color = 2'b00;
		14'h3120: color = 2'b00;
		14'h3121: color = 2'b00;
		14'h3122: color = 2'b00;
		14'h3123: color = 2'b00;
		14'h3124: color = 2'b00;
		14'h3125: color = 2'b00;
		14'h3126: color = 2'b01;
		14'h3127: color = 2'b00;
		14'h3128: color = 2'b00;
		14'h3129: color = 2'b01;
		14'h312a: color = 2'b01;
		14'h312b: color = 2'b00;
		14'h312c: color = 2'b00;
		14'h312d: color = 2'b00;
		14'h312e: color = 2'b00;
		14'h312f: color = 2'b00;
		14'h3130: color = 2'b00;
		14'h3131: color = 2'b01;
		14'h3132: color = 2'b11;
		14'h3133: color = 2'b11;
		14'h3134: color = 2'b11;
		14'h3135: color = 2'b11;
		14'h3136: color = 2'b11;
		14'h3137: color = 2'b11;
		14'h3138: color = 2'b11;
		14'h3139: color = 2'b11;
		14'h313a: color = 2'b11;
		14'h313b: color = 2'b10;
		14'h313c: color = 2'b01;
		14'h313d: color = 2'b10;
		14'h313e: color = 2'b01;
		14'h313f: color = 2'b01;
		14'h3140: color = 2'b01;
		14'h3141: color = 2'b01;
		14'h3142: color = 2'b01;
		14'h3143: color = 2'b01;
		14'h3144: color = 2'b01;
		14'h3145: color = 2'b01;
		14'h3146: color = 2'b00;
		14'h3147: color = 2'b00;
		14'h3148: color = 2'b00;
		14'h3149: color = 2'b00;
		14'h314a: color = 2'b00;
		14'h314b: color = 2'b00;
		14'h314c: color = 2'b00;
		14'h314d: color = 2'b00;
		14'h314e: color = 2'b10;
		14'h314f: color = 2'b10;
		14'h3150: color = 2'b11;
		14'h3151: color = 2'b01;
		14'h3152: color = 2'b00;
		14'h3153: color = 2'b00;
		14'h3154: color = 2'b00;
		14'h3155: color = 2'b00;
		14'h3156: color = 2'b00;
		14'h3157: color = 2'b00;
		14'h3158: color = 2'b00;
		14'h3159: color = 2'b00;
		14'h315a: color = 2'b00;
		14'h315b: color = 2'b00;
		14'h315c: color = 2'b00;
		14'h315d: color = 2'b00;
		14'h315e: color = 2'b00;
		14'h315f: color = 2'b00;
		14'h3160: color = 2'b00;
		14'h3161: color = 2'b00;
		14'h3162: color = 2'b00;
		14'h3163: color = 2'b00;
		14'h3164: color = 2'b00;
		14'h3165: color = 2'b00;
		14'h3166: color = 2'b00;
		14'h3167: color = 2'b00;
		14'h3168: color = 2'b00;
		14'h3169: color = 2'b00;
		14'h316a: color = 2'b00;
		14'h316b: color = 2'b00;
		14'h316c: color = 2'b00;
		14'h316d: color = 2'b00;
		14'h316e: color = 2'b00;
		14'h316f: color = 2'b00;
		14'h3170: color = 2'b00;
		14'h3171: color = 2'b10;
		14'h3172: color = 2'b11;
		14'h3173: color = 2'b11;
		14'h3174: color = 2'b11;
		14'h3175: color = 2'b11;
		14'h3176: color = 2'b11;
		14'h3177: color = 2'b11;
		14'h3178: color = 2'b11;
		14'h3179: color = 2'b11;
		14'h317a: color = 2'b11;
		14'h317b: color = 2'b11;
		14'h317c: color = 2'b11;
		14'h317d: color = 2'b11;
		14'h317e: color = 2'b11;
		14'h317f: color = 2'b11;
		14'h3180: color = 2'b01;
		14'h3181: color = 2'b01;
		14'h3182: color = 2'b00;
		14'h3183: color = 2'b00;
		14'h3184: color = 2'b01;
		14'h3185: color = 2'b00;
		14'h3186: color = 2'b00;
		14'h3187: color = 2'b00;
		14'h3188: color = 2'b00;
		14'h3189: color = 2'b00;
		14'h318a: color = 2'b00;
		14'h318b: color = 2'b00;
		14'h318c: color = 2'b00;
		14'h318d: color = 2'b00;
		14'h318e: color = 2'b00;
		14'h318f: color = 2'b00;
		14'h3190: color = 2'b00;
		14'h3191: color = 2'b00;
		14'h3192: color = 2'b00;
		14'h3193: color = 2'b00;
		14'h3194: color = 2'b00;
		14'h3195: color = 2'b00;
		14'h3196: color = 2'b00;
		14'h3197: color = 2'b00;
		14'h3198: color = 2'b00;
		14'h3199: color = 2'b00;
		14'h319a: color = 2'b00;
		14'h319b: color = 2'b00;
		14'h319c: color = 2'b00;
		14'h319d: color = 2'b00;
		14'h319e: color = 2'b00;
		14'h319f: color = 2'b00;
		14'h31a0: color = 2'b00;
		14'h31a1: color = 2'b00;
		14'h31a2: color = 2'b00;
		14'h31a3: color = 2'b00;
		14'h31a4: color = 2'b00;
		14'h31a5: color = 2'b00;
		14'h31a6: color = 2'b00;
		14'h31a7: color = 2'b00;
		14'h31a8: color = 2'b00;
		14'h31a9: color = 2'b01;
		14'h31aa: color = 2'b00;
		14'h31ab: color = 2'b00;
		14'h31ac: color = 2'b00;
		14'h31ad: color = 2'b00;
		14'h31ae: color = 2'b00;
		14'h31af: color = 2'b00;
		14'h31b0: color = 2'b00;
		14'h31b1: color = 2'b00;
		14'h31b2: color = 2'b10;
		14'h31b3: color = 2'b11;
		14'h31b4: color = 2'b11;
		14'h31b5: color = 2'b11;
		14'h31b6: color = 2'b11;
		14'h31b7: color = 2'b11;
		14'h31b8: color = 2'b11;
		14'h31b9: color = 2'b11;
		14'h31ba: color = 2'b11;
		14'h31bb: color = 2'b11;
		14'h31bc: color = 2'b10;
		14'h31bd: color = 2'b10;
		14'h31be: color = 2'b01;
		14'h31bf: color = 2'b01;
		14'h31c0: color = 2'b01;
		14'h31c1: color = 2'b01;
		14'h31c2: color = 2'b10;
		14'h31c3: color = 2'b01;
		14'h31c4: color = 2'b01;
		14'h31c5: color = 2'b01;
		14'h31c6: color = 2'b01;
		14'h31c7: color = 2'b00;
		14'h31c8: color = 2'b00;
		14'h31c9: color = 2'b00;
		14'h31ca: color = 2'b00;
		14'h31cb: color = 2'b00;
		14'h31cc: color = 2'b00;
		14'h31cd: color = 2'b01;
		14'h31ce: color = 2'b10;
		14'h31cf: color = 2'b11;
		14'h31d0: color = 2'b11;
		14'h31d1: color = 2'b01;
		14'h31d2: color = 2'b00;
		14'h31d3: color = 2'b00;
		14'h31d4: color = 2'b00;
		14'h31d5: color = 2'b00;
		14'h31d6: color = 2'b00;
		14'h31d7: color = 2'b00;
		14'h31d8: color = 2'b00;
		14'h31d9: color = 2'b00;
		14'h31da: color = 2'b00;
		14'h31db: color = 2'b00;
		14'h31dc: color = 2'b00;
		14'h31dd: color = 2'b00;
		14'h31de: color = 2'b00;
		14'h31df: color = 2'b00;
		14'h31e0: color = 2'b00;
		14'h31e1: color = 2'b00;
		14'h31e2: color = 2'b00;
		14'h31e3: color = 2'b00;
		14'h31e4: color = 2'b00;
		14'h31e5: color = 2'b00;
		14'h31e6: color = 2'b00;
		14'h31e7: color = 2'b00;
		14'h31e8: color = 2'b00;
		14'h31e9: color = 2'b00;
		14'h31ea: color = 2'b00;
		14'h31eb: color = 2'b00;
		14'h31ec: color = 2'b00;
		14'h31ed: color = 2'b00;
		14'h31ee: color = 2'b00;
		14'h31ef: color = 2'b00;
		14'h31f0: color = 2'b00;
		14'h31f1: color = 2'b00;
		14'h31f2: color = 2'b00;
		14'h31f3: color = 2'b11;
		14'h31f4: color = 2'b11;
		14'h31f5: color = 2'b11;
		14'h31f6: color = 2'b11;
		14'h31f7: color = 2'b11;
		14'h31f8: color = 2'b11;
		14'h31f9: color = 2'b11;
		14'h31fa: color = 2'b11;
		14'h31fb: color = 2'b11;
		14'h31fc: color = 2'b11;
		14'h31fd: color = 2'b11;
		14'h31fe: color = 2'b11;
		14'h31ff: color = 2'b11;
		14'h3200: color = 2'b00;
		14'h3201: color = 2'b00;
		14'h3202: color = 2'b01;
		14'h3203: color = 2'b00;
		14'h3204: color = 2'b00;
		14'h3205: color = 2'b01;
		14'h3206: color = 2'b00;
		14'h3207: color = 2'b01;
		14'h3208: color = 2'b01;
		14'h3209: color = 2'b00;
		14'h320a: color = 2'b00;
		14'h320b: color = 2'b01;
		14'h320c: color = 2'b00;
		14'h320d: color = 2'b00;
		14'h320e: color = 2'b00;
		14'h320f: color = 2'b00;
		14'h3210: color = 2'b00;
		14'h3211: color = 2'b00;
		14'h3212: color = 2'b00;
		14'h3213: color = 2'b00;
		14'h3214: color = 2'b00;
		14'h3215: color = 2'b00;
		14'h3216: color = 2'b00;
		14'h3217: color = 2'b00;
		14'h3218: color = 2'b00;
		14'h3219: color = 2'b00;
		14'h321a: color = 2'b00;
		14'h321b: color = 2'b00;
		14'h321c: color = 2'b00;
		14'h321d: color = 2'b00;
		14'h321e: color = 2'b00;
		14'h321f: color = 2'b00;
		14'h3220: color = 2'b00;
		14'h3221: color = 2'b00;
		14'h3222: color = 2'b00;
		14'h3223: color = 2'b00;
		14'h3224: color = 2'b00;
		14'h3225: color = 2'b00;
		14'h3226: color = 2'b00;
		14'h3227: color = 2'b01;
		14'h3228: color = 2'b01;
		14'h3229: color = 2'b00;
		14'h322a: color = 2'b00;
		14'h322b: color = 2'b00;
		14'h322c: color = 2'b00;
		14'h322d: color = 2'b00;
		14'h322e: color = 2'b00;
		14'h322f: color = 2'b00;
		14'h3230: color = 2'b00;
		14'h3231: color = 2'b00;
		14'h3232: color = 2'b01;
		14'h3233: color = 2'b11;
		14'h3234: color = 2'b11;
		14'h3235: color = 2'b11;
		14'h3236: color = 2'b11;
		14'h3237: color = 2'b11;
		14'h3238: color = 2'b11;
		14'h3239: color = 2'b11;
		14'h323a: color = 2'b11;
		14'h323b: color = 2'b11;
		14'h323c: color = 2'b11;
		14'h323d: color = 2'b10;
		14'h323e: color = 2'b01;
		14'h323f: color = 2'b01;
		14'h3240: color = 2'b01;
		14'h3241: color = 2'b01;
		14'h3242: color = 2'b01;
		14'h3243: color = 2'b01;
		14'h3244: color = 2'b01;
		14'h3245: color = 2'b01;
		14'h3246: color = 2'b00;
		14'h3247: color = 2'b00;
		14'h3248: color = 2'b00;
		14'h3249: color = 2'b00;
		14'h324a: color = 2'b00;
		14'h324b: color = 2'b01;
		14'h324c: color = 2'b01;
		14'h324d: color = 2'b10;
		14'h324e: color = 2'b11;
		14'h324f: color = 2'b11;
		14'h3250: color = 2'b10;
		14'h3251: color = 2'b10;
		14'h3252: color = 2'b00;
		14'h3253: color = 2'b00;
		14'h3254: color = 2'b00;
		14'h3255: color = 2'b00;
		14'h3256: color = 2'b00;
		14'h3257: color = 2'b00;
		14'h3258: color = 2'b00;
		14'h3259: color = 2'b00;
		14'h325a: color = 2'b00;
		14'h325b: color = 2'b00;
		14'h325c: color = 2'b00;
		14'h325d: color = 2'b00;
		14'h325e: color = 2'b00;
		14'h325f: color = 2'b00;
		14'h3260: color = 2'b00;
		14'h3261: color = 2'b00;
		14'h3262: color = 2'b00;
		14'h3263: color = 2'b00;
		14'h3264: color = 2'b00;
		14'h3265: color = 2'b00;
		14'h3266: color = 2'b00;
		14'h3267: color = 2'b00;
		14'h3268: color = 2'b00;
		14'h3269: color = 2'b00;
		14'h326a: color = 2'b00;
		14'h326b: color = 2'b00;
		14'h326c: color = 2'b00;
		14'h326d: color = 2'b00;
		14'h326e: color = 2'b00;
		14'h326f: color = 2'b00;
		14'h3270: color = 2'b00;
		14'h3271: color = 2'b00;
		14'h3272: color = 2'b00;
		14'h3273: color = 2'b01;
		14'h3274: color = 2'b11;
		14'h3275: color = 2'b11;
		14'h3276: color = 2'b11;
		14'h3277: color = 2'b11;
		14'h3278: color = 2'b11;
		14'h3279: color = 2'b11;
		14'h327a: color = 2'b11;
		14'h327b: color = 2'b11;
		14'h327c: color = 2'b11;
		14'h327d: color = 2'b11;
		14'h327e: color = 2'b11;
		14'h327f: color = 2'b11;
		14'h3280: color = 2'b00;
		14'h3281: color = 2'b00;
		14'h3282: color = 2'b01;
		14'h3283: color = 2'b00;
		14'h3284: color = 2'b00;
		14'h3285: color = 2'b01;
		14'h3286: color = 2'b00;
		14'h3287: color = 2'b00;
		14'h3288: color = 2'b00;
		14'h3289: color = 2'b01;
		14'h328a: color = 2'b00;
		14'h328b: color = 2'b00;
		14'h328c: color = 2'b00;
		14'h328d: color = 2'b00;
		14'h328e: color = 2'b00;
		14'h328f: color = 2'b00;
		14'h3290: color = 2'b00;
		14'h3291: color = 2'b00;
		14'h3292: color = 2'b00;
		14'h3293: color = 2'b00;
		14'h3294: color = 2'b00;
		14'h3295: color = 2'b00;
		14'h3296: color = 2'b00;
		14'h3297: color = 2'b00;
		14'h3298: color = 2'b00;
		14'h3299: color = 2'b00;
		14'h329a: color = 2'b00;
		14'h329b: color = 2'b00;
		14'h329c: color = 2'b00;
		14'h329d: color = 2'b00;
		14'h329e: color = 2'b00;
		14'h329f: color = 2'b00;
		14'h32a0: color = 2'b00;
		14'h32a1: color = 2'b00;
		14'h32a2: color = 2'b00;
		14'h32a3: color = 2'b00;
		14'h32a4: color = 2'b00;
		14'h32a5: color = 2'b00;
		14'h32a6: color = 2'b01;
		14'h32a7: color = 2'b00;
		14'h32a8: color = 2'b00;
		14'h32a9: color = 2'b01;
		14'h32aa: color = 2'b00;
		14'h32ab: color = 2'b00;
		14'h32ac: color = 2'b00;
		14'h32ad: color = 2'b00;
		14'h32ae: color = 2'b00;
		14'h32af: color = 2'b00;
		14'h32b0: color = 2'b00;
		14'h32b1: color = 2'b00;
		14'h32b2: color = 2'b01;
		14'h32b3: color = 2'b10;
		14'h32b4: color = 2'b11;
		14'h32b5: color = 2'b11;
		14'h32b6: color = 2'b11;
		14'h32b7: color = 2'b11;
		14'h32b8: color = 2'b11;
		14'h32b9: color = 2'b11;
		14'h32ba: color = 2'b10;
		14'h32bb: color = 2'b11;
		14'h32bc: color = 2'b11;
		14'h32bd: color = 2'b10;
		14'h32be: color = 2'b10;
		14'h32bf: color = 2'b01;
		14'h32c0: color = 2'b01;
		14'h32c1: color = 2'b00;
		14'h32c2: color = 2'b01;
		14'h32c3: color = 2'b01;
		14'h32c4: color = 2'b01;
		14'h32c5: color = 2'b01;
		14'h32c6: color = 2'b00;
		14'h32c7: color = 2'b01;
		14'h32c8: color = 2'b01;
		14'h32c9: color = 2'b00;
		14'h32ca: color = 2'b01;
		14'h32cb: color = 2'b01;
		14'h32cc: color = 2'b10;
		14'h32cd: color = 2'b11;
		14'h32ce: color = 2'b11;
		14'h32cf: color = 2'b10;
		14'h32d0: color = 2'b11;
		14'h32d1: color = 2'b10;
		14'h32d2: color = 2'b00;
		14'h32d3: color = 2'b00;
		14'h32d4: color = 2'b00;
		14'h32d5: color = 2'b00;
		14'h32d6: color = 2'b00;
		14'h32d7: color = 2'b00;
		14'h32d8: color = 2'b00;
		14'h32d9: color = 2'b00;
		14'h32da: color = 2'b00;
		14'h32db: color = 2'b00;
		14'h32dc: color = 2'b00;
		14'h32dd: color = 2'b00;
		14'h32de: color = 2'b00;
		14'h32df: color = 2'b00;
		14'h32e0: color = 2'b00;
		14'h32e1: color = 2'b00;
		14'h32e2: color = 2'b00;
		14'h32e3: color = 2'b00;
		14'h32e4: color = 2'b00;
		14'h32e5: color = 2'b00;
		14'h32e6: color = 2'b00;
		14'h32e7: color = 2'b00;
		14'h32e8: color = 2'b00;
		14'h32e9: color = 2'b00;
		14'h32ea: color = 2'b00;
		14'h32eb: color = 2'b00;
		14'h32ec: color = 2'b00;
		14'h32ed: color = 2'b00;
		14'h32ee: color = 2'b00;
		14'h32ef: color = 2'b00;
		14'h32f0: color = 2'b00;
		14'h32f1: color = 2'b00;
		14'h32f2: color = 2'b00;
		14'h32f3: color = 2'b00;
		14'h32f4: color = 2'b00;
		14'h32f5: color = 2'b11;
		14'h32f6: color = 2'b11;
		14'h32f7: color = 2'b11;
		14'h32f8: color = 2'b11;
		14'h32f9: color = 2'b11;
		14'h32fa: color = 2'b11;
		14'h32fb: color = 2'b11;
		14'h32fc: color = 2'b11;
		14'h32fd: color = 2'b11;
		14'h32fe: color = 2'b11;
		14'h32ff: color = 2'b11;
		14'h3300: color = 2'b01;
		14'h3301: color = 2'b00;
		14'h3302: color = 2'b00;
		14'h3303: color = 2'b01;
		14'h3304: color = 2'b00;
		14'h3305: color = 2'b00;
		14'h3306: color = 2'b00;
		14'h3307: color = 2'b00;
		14'h3308: color = 2'b00;
		14'h3309: color = 2'b00;
		14'h330a: color = 2'b00;
		14'h330b: color = 2'b00;
		14'h330c: color = 2'b00;
		14'h330d: color = 2'b00;
		14'h330e: color = 2'b01;
		14'h330f: color = 2'b00;
		14'h3310: color = 2'b00;
		14'h3311: color = 2'b00;
		14'h3312: color = 2'b00;
		14'h3313: color = 2'b00;
		14'h3314: color = 2'b00;
		14'h3315: color = 2'b00;
		14'h3316: color = 2'b00;
		14'h3317: color = 2'b00;
		14'h3318: color = 2'b00;
		14'h3319: color = 2'b00;
		14'h331a: color = 2'b00;
		14'h331b: color = 2'b00;
		14'h331c: color = 2'b00;
		14'h331d: color = 2'b00;
		14'h331e: color = 2'b00;
		14'h331f: color = 2'b00;
		14'h3320: color = 2'b00;
		14'h3321: color = 2'b00;
		14'h3322: color = 2'b00;
		14'h3323: color = 2'b00;
		14'h3324: color = 2'b00;
		14'h3325: color = 2'b00;
		14'h3326: color = 2'b00;
		14'h3327: color = 2'b00;
		14'h3328: color = 2'b00;
		14'h3329: color = 2'b00;
		14'h332a: color = 2'b00;
		14'h332b: color = 2'b00;
		14'h332c: color = 2'b00;
		14'h332d: color = 2'b00;
		14'h332e: color = 2'b00;
		14'h332f: color = 2'b00;
		14'h3330: color = 2'b00;
		14'h3331: color = 2'b00;
		14'h3332: color = 2'b00;
		14'h3333: color = 2'b01;
		14'h3334: color = 2'b11;
		14'h3335: color = 2'b11;
		14'h3336: color = 2'b11;
		14'h3337: color = 2'b11;
		14'h3338: color = 2'b11;
		14'h3339: color = 2'b11;
		14'h333a: color = 2'b11;
		14'h333b: color = 2'b10;
		14'h333c: color = 2'b10;
		14'h333d: color = 2'b11;
		14'h333e: color = 2'b10;
		14'h333f: color = 2'b01;
		14'h3340: color = 2'b00;
		14'h3341: color = 2'b01;
		14'h3342: color = 2'b00;
		14'h3343: color = 2'b01;
		14'h3344: color = 2'b01;
		14'h3345: color = 2'b01;
		14'h3346: color = 2'b01;
		14'h3347: color = 2'b00;
		14'h3348: color = 2'b00;
		14'h3349: color = 2'b01;
		14'h334a: color = 2'b01;
		14'h334b: color = 2'b10;
		14'h334c: color = 2'b11;
		14'h334d: color = 2'b11;
		14'h334e: color = 2'b10;
		14'h334f: color = 2'b11;
		14'h3350: color = 2'b10;
		14'h3351: color = 2'b10;
		14'h3352: color = 2'b00;
		14'h3353: color = 2'b00;
		14'h3354: color = 2'b00;
		14'h3355: color = 2'b00;
		14'h3356: color = 2'b00;
		14'h3357: color = 2'b00;
		14'h3358: color = 2'b00;
		14'h3359: color = 2'b00;
		14'h335a: color = 2'b00;
		14'h335b: color = 2'b00;
		14'h335c: color = 2'b00;
		14'h335d: color = 2'b00;
		14'h335e: color = 2'b00;
		14'h335f: color = 2'b00;
		14'h3360: color = 2'b00;
		14'h3361: color = 2'b00;
		14'h3362: color = 2'b00;
		14'h3363: color = 2'b00;
		14'h3364: color = 2'b00;
		14'h3365: color = 2'b00;
		14'h3366: color = 2'b00;
		14'h3367: color = 2'b00;
		14'h3368: color = 2'b00;
		14'h3369: color = 2'b00;
		14'h336a: color = 2'b00;
		14'h336b: color = 2'b00;
		14'h336c: color = 2'b00;
		14'h336d: color = 2'b00;
		14'h336e: color = 2'b00;
		14'h336f: color = 2'b00;
		14'h3370: color = 2'b00;
		14'h3371: color = 2'b00;
		14'h3372: color = 2'b00;
		14'h3373: color = 2'b00;
		14'h3374: color = 2'b00;
		14'h3375: color = 2'b10;
		14'h3376: color = 2'b11;
		14'h3377: color = 2'b11;
		14'h3378: color = 2'b11;
		14'h3379: color = 2'b11;
		14'h337a: color = 2'b11;
		14'h337b: color = 2'b11;
		14'h337c: color = 2'b11;
		14'h337d: color = 2'b11;
		14'h337e: color = 2'b11;
		14'h337f: color = 2'b11;
		14'h3380: color = 2'b00;
		14'h3381: color = 2'b00;
		14'h3382: color = 2'b00;
		14'h3383: color = 2'b01;
		14'h3384: color = 2'b00;
		14'h3385: color = 2'b00;
		14'h3386: color = 2'b01;
		14'h3387: color = 2'b00;
		14'h3388: color = 2'b00;
		14'h3389: color = 2'b01;
		14'h338a: color = 2'b00;
		14'h338b: color = 2'b00;
		14'h338c: color = 2'b01;
		14'h338d: color = 2'b00;
		14'h338e: color = 2'b00;
		14'h338f: color = 2'b00;
		14'h3390: color = 2'b00;
		14'h3391: color = 2'b00;
		14'h3392: color = 2'b00;
		14'h3393: color = 2'b00;
		14'h3394: color = 2'b00;
		14'h3395: color = 2'b00;
		14'h3396: color = 2'b00;
		14'h3397: color = 2'b00;
		14'h3398: color = 2'b00;
		14'h3399: color = 2'b00;
		14'h339a: color = 2'b00;
		14'h339b: color = 2'b00;
		14'h339c: color = 2'b00;
		14'h339d: color = 2'b00;
		14'h339e: color = 2'b00;
		14'h339f: color = 2'b00;
		14'h33a0: color = 2'b00;
		14'h33a1: color = 2'b00;
		14'h33a2: color = 2'b00;
		14'h33a3: color = 2'b00;
		14'h33a4: color = 2'b00;
		14'h33a5: color = 2'b00;
		14'h33a6: color = 2'b00;
		14'h33a7: color = 2'b00;
		14'h33a8: color = 2'b00;
		14'h33a9: color = 2'b00;
		14'h33aa: color = 2'b00;
		14'h33ab: color = 2'b00;
		14'h33ac: color = 2'b00;
		14'h33ad: color = 2'b00;
		14'h33ae: color = 2'b00;
		14'h33af: color = 2'b00;
		14'h33b0: color = 2'b00;
		14'h33b1: color = 2'b00;
		14'h33b2: color = 2'b00;
		14'h33b3: color = 2'b01;
		14'h33b4: color = 2'b10;
		14'h33b5: color = 2'b11;
		14'h33b6: color = 2'b11;
		14'h33b7: color = 2'b11;
		14'h33b8: color = 2'b11;
		14'h33b9: color = 2'b11;
		14'h33ba: color = 2'b11;
		14'h33bb: color = 2'b11;
		14'h33bc: color = 2'b10;
		14'h33bd: color = 2'b10;
		14'h33be: color = 2'b11;
		14'h33bf: color = 2'b10;
		14'h33c0: color = 2'b10;
		14'h33c1: color = 2'b00;
		14'h33c2: color = 2'b01;
		14'h33c3: color = 2'b01;
		14'h33c4: color = 2'b00;
		14'h33c5: color = 2'b01;
		14'h33c6: color = 2'b00;
		14'h33c7: color = 2'b01;
		14'h33c8: color = 2'b01;
		14'h33c9: color = 2'b01;
		14'h33ca: color = 2'b10;
		14'h33cb: color = 2'b11;
		14'h33cc: color = 2'b10;
		14'h33cd: color = 2'b11;
		14'h33ce: color = 2'b11;
		14'h33cf: color = 2'b10;
		14'h33d0: color = 2'b11;
		14'h33d1: color = 2'b10;
		14'h33d2: color = 2'b00;
		14'h33d3: color = 2'b00;
		14'h33d4: color = 2'b00;
		14'h33d5: color = 2'b00;
		14'h33d6: color = 2'b00;
		14'h33d7: color = 2'b00;
		14'h33d8: color = 2'b00;
		14'h33d9: color = 2'b00;
		14'h33da: color = 2'b00;
		14'h33db: color = 2'b00;
		14'h33dc: color = 2'b00;
		14'h33dd: color = 2'b00;
		14'h33de: color = 2'b00;
		14'h33df: color = 2'b00;
		14'h33e0: color = 2'b00;
		14'h33e1: color = 2'b00;
		14'h33e2: color = 2'b00;
		14'h33e3: color = 2'b00;
		14'h33e4: color = 2'b00;
		14'h33e5: color = 2'b00;
		14'h33e6: color = 2'b00;
		14'h33e7: color = 2'b00;
		14'h33e8: color = 2'b00;
		14'h33e9: color = 2'b00;
		14'h33ea: color = 2'b00;
		14'h33eb: color = 2'b00;
		14'h33ec: color = 2'b00;
		14'h33ed: color = 2'b00;
		14'h33ee: color = 2'b00;
		14'h33ef: color = 2'b00;
		14'h33f0: color = 2'b00;
		14'h33f1: color = 2'b00;
		14'h33f2: color = 2'b00;
		14'h33f3: color = 2'b00;
		14'h33f4: color = 2'b00;
		14'h33f5: color = 2'b00;
		14'h33f6: color = 2'b11;
		14'h33f7: color = 2'b11;
		14'h33f8: color = 2'b11;
		14'h33f9: color = 2'b11;
		14'h33fa: color = 2'b11;
		14'h33fb: color = 2'b11;
		14'h33fc: color = 2'b11;
		14'h33fd: color = 2'b11;
		14'h33fe: color = 2'b11;
		14'h33ff: color = 2'b11;
		14'h3400: color = 2'b00;
		14'h3401: color = 2'b00;
		14'h3402: color = 2'b00;
		14'h3403: color = 2'b01;
		14'h3404: color = 2'b00;
		14'h3405: color = 2'b00;
		14'h3406: color = 2'b01;
		14'h3407: color = 2'b00;
		14'h3408: color = 2'b00;
		14'h3409: color = 2'b01;
		14'h340a: color = 2'b00;
		14'h340b: color = 2'b00;
		14'h340c: color = 2'b01;
		14'h340d: color = 2'b00;
		14'h340e: color = 2'b00;
		14'h340f: color = 2'b00;
		14'h3410: color = 2'b00;
		14'h3411: color = 2'b00;
		14'h3412: color = 2'b00;
		14'h3413: color = 2'b00;
		14'h3414: color = 2'b00;
		14'h3415: color = 2'b00;
		14'h3416: color = 2'b00;
		14'h3417: color = 2'b00;
		14'h3418: color = 2'b00;
		14'h3419: color = 2'b00;
		14'h341a: color = 2'b00;
		14'h341b: color = 2'b00;
		14'h341c: color = 2'b00;
		14'h341d: color = 2'b00;
		14'h341e: color = 2'b00;
		14'h341f: color = 2'b00;
		14'h3420: color = 2'b00;
		14'h3421: color = 2'b00;
		14'h3422: color = 2'b00;
		14'h3423: color = 2'b00;
		14'h3424: color = 2'b00;
		14'h3425: color = 2'b00;
		14'h3426: color = 2'b00;
		14'h3427: color = 2'b00;
		14'h3428: color = 2'b00;
		14'h3429: color = 2'b00;
		14'h342a: color = 2'b00;
		14'h342b: color = 2'b00;
		14'h342c: color = 2'b00;
		14'h342d: color = 2'b00;
		14'h342e: color = 2'b00;
		14'h342f: color = 2'b00;
		14'h3430: color = 2'b00;
		14'h3431: color = 2'b00;
		14'h3432: color = 2'b00;
		14'h3433: color = 2'b01;
		14'h3434: color = 2'b10;
		14'h3435: color = 2'b11;
		14'h3436: color = 2'b11;
		14'h3437: color = 2'b11;
		14'h3438: color = 2'b11;
		14'h3439: color = 2'b11;
		14'h343a: color = 2'b11;
		14'h343b: color = 2'b11;
		14'h343c: color = 2'b10;
		14'h343d: color = 2'b10;
		14'h343e: color = 2'b11;
		14'h343f: color = 2'b10;
		14'h3440: color = 2'b10;
		14'h3441: color = 2'b00;
		14'h3442: color = 2'b01;
		14'h3443: color = 2'b01;
		14'h3444: color = 2'b00;
		14'h3445: color = 2'b01;
		14'h3446: color = 2'b00;
		14'h3447: color = 2'b01;
		14'h3448: color = 2'b01;
		14'h3449: color = 2'b01;
		14'h344a: color = 2'b10;
		14'h344b: color = 2'b11;
		14'h344c: color = 2'b10;
		14'h344d: color = 2'b11;
		14'h344e: color = 2'b11;
		14'h344f: color = 2'b10;
		14'h3450: color = 2'b11;
		14'h3451: color = 2'b10;
		14'h3452: color = 2'b00;
		14'h3453: color = 2'b00;
		14'h3454: color = 2'b00;
		14'h3455: color = 2'b00;
		14'h3456: color = 2'b00;
		14'h3457: color = 2'b00;
		14'h3458: color = 2'b00;
		14'h3459: color = 2'b00;
		14'h345a: color = 2'b00;
		14'h345b: color = 2'b00;
		14'h345c: color = 2'b00;
		14'h345d: color = 2'b00;
		14'h345e: color = 2'b00;
		14'h345f: color = 2'b00;
		14'h3460: color = 2'b00;
		14'h3461: color = 2'b00;
		14'h3462: color = 2'b00;
		14'h3463: color = 2'b00;
		14'h3464: color = 2'b00;
		14'h3465: color = 2'b00;
		14'h3466: color = 2'b00;
		14'h3467: color = 2'b00;
		14'h3468: color = 2'b00;
		14'h3469: color = 2'b00;
		14'h346a: color = 2'b00;
		14'h346b: color = 2'b00;
		14'h346c: color = 2'b00;
		14'h346d: color = 2'b00;
		14'h346e: color = 2'b00;
		14'h346f: color = 2'b00;
		14'h3470: color = 2'b00;
		14'h3471: color = 2'b00;
		14'h3472: color = 2'b00;
		14'h3473: color = 2'b00;
		14'h3474: color = 2'b00;
		14'h3475: color = 2'b00;
		14'h3476: color = 2'b11;
		14'h3477: color = 2'b11;
		14'h3478: color = 2'b11;
		14'h3479: color = 2'b11;
		14'h347a: color = 2'b11;
		14'h347b: color = 2'b11;
		14'h347c: color = 2'b11;
		14'h347d: color = 2'b11;
		14'h347e: color = 2'b11;
		14'h347f: color = 2'b11;
		14'h3480: color = 2'b00;
		14'h3481: color = 2'b01;
		14'h3482: color = 2'b00;
		14'h3483: color = 2'b00;
		14'h3484: color = 2'b00;
		14'h3485: color = 2'b00;
		14'h3486: color = 2'b00;
		14'h3487: color = 2'b00;
		14'h3488: color = 2'b00;
		14'h3489: color = 2'b00;
		14'h348a: color = 2'b00;
		14'h348b: color = 2'b00;
		14'h348c: color = 2'b00;
		14'h348d: color = 2'b00;
		14'h348e: color = 2'b00;
		14'h348f: color = 2'b00;
		14'h3490: color = 2'b00;
		14'h3491: color = 2'b00;
		14'h3492: color = 2'b00;
		14'h3493: color = 2'b00;
		14'h3494: color = 2'b00;
		14'h3495: color = 2'b00;
		14'h3496: color = 2'b00;
		14'h3497: color = 2'b00;
		14'h3498: color = 2'b00;
		14'h3499: color = 2'b00;
		14'h349a: color = 2'b00;
		14'h349b: color = 2'b00;
		14'h349c: color = 2'b00;
		14'h349d: color = 2'b00;
		14'h349e: color = 2'b00;
		14'h349f: color = 2'b00;
		14'h34a0: color = 2'b00;
		14'h34a1: color = 2'b00;
		14'h34a2: color = 2'b00;
		14'h34a3: color = 2'b00;
		14'h34a4: color = 2'b00;
		14'h34a5: color = 2'b00;
		14'h34a6: color = 2'b00;
		14'h34a7: color = 2'b00;
		14'h34a8: color = 2'b00;
		14'h34a9: color = 2'b00;
		14'h34aa: color = 2'b00;
		14'h34ab: color = 2'b00;
		14'h34ac: color = 2'b00;
		14'h34ad: color = 2'b00;
		14'h34ae: color = 2'b00;
		14'h34af: color = 2'b00;
		14'h34b0: color = 2'b00;
		14'h34b1: color = 2'b00;
		14'h34b2: color = 2'b00;
		14'h34b3: color = 2'b00;
		14'h34b4: color = 2'b01;
		14'h34b5: color = 2'b10;
		14'h34b6: color = 2'b11;
		14'h34b7: color = 2'b11;
		14'h34b8: color = 2'b11;
		14'h34b9: color = 2'b11;
		14'h34ba: color = 2'b11;
		14'h34bb: color = 2'b10;
		14'h34bc: color = 2'b11;
		14'h34bd: color = 2'b10;
		14'h34be: color = 2'b10;
		14'h34bf: color = 2'b11;
		14'h34c0: color = 2'b11;
		14'h34c1: color = 2'b10;
		14'h34c2: color = 2'b01;
		14'h34c3: color = 2'b01;
		14'h34c4: color = 2'b00;
		14'h34c5: color = 2'b01;
		14'h34c6: color = 2'b01;
		14'h34c7: color = 2'b10;
		14'h34c8: color = 2'b10;
		14'h34c9: color = 2'b11;
		14'h34ca: color = 2'b11;
		14'h34cb: color = 2'b11;
		14'h34cc: color = 2'b11;
		14'h34cd: color = 2'b10;
		14'h34ce: color = 2'b11;
		14'h34cf: color = 2'b11;
		14'h34d0: color = 2'b10;
		14'h34d1: color = 2'b11;
		14'h34d2: color = 2'b00;
		14'h34d3: color = 2'b00;
		14'h34d4: color = 2'b00;
		14'h34d5: color = 2'b00;
		14'h34d6: color = 2'b00;
		14'h34d7: color = 2'b00;
		14'h34d8: color = 2'b00;
		14'h34d9: color = 2'b00;
		14'h34da: color = 2'b00;
		14'h34db: color = 2'b00;
		14'h34dc: color = 2'b00;
		14'h34dd: color = 2'b00;
		14'h34de: color = 2'b00;
		14'h34df: color = 2'b00;
		14'h34e0: color = 2'b00;
		14'h34e1: color = 2'b00;
		14'h34e2: color = 2'b00;
		14'h34e3: color = 2'b00;
		14'h34e4: color = 2'b00;
		14'h34e5: color = 2'b00;
		14'h34e6: color = 2'b00;
		14'h34e7: color = 2'b00;
		14'h34e8: color = 2'b00;
		14'h34e9: color = 2'b00;
		14'h34ea: color = 2'b00;
		14'h34eb: color = 2'b00;
		14'h34ec: color = 2'b00;
		14'h34ed: color = 2'b00;
		14'h34ee: color = 2'b00;
		14'h34ef: color = 2'b00;
		14'h34f0: color = 2'b00;
		14'h34f1: color = 2'b00;
		14'h34f2: color = 2'b00;
		14'h34f3: color = 2'b00;
		14'h34f4: color = 2'b00;
		14'h34f5: color = 2'b00;
		14'h34f6: color = 2'b10;
		14'h34f7: color = 2'b11;
		14'h34f8: color = 2'b11;
		14'h34f9: color = 2'b11;
		14'h34fa: color = 2'b11;
		14'h34fb: color = 2'b11;
		14'h34fc: color = 2'b11;
		14'h34fd: color = 2'b11;
		14'h34fe: color = 2'b11;
		14'h34ff: color = 2'b11;
		14'h3500: color = 2'b00;
		14'h3501: color = 2'b01;
		14'h3502: color = 2'b00;
		14'h3503: color = 2'b01;
		14'h3504: color = 2'b00;
		14'h3505: color = 2'b00;
		14'h3506: color = 2'b01;
		14'h3507: color = 2'b00;
		14'h3508: color = 2'b00;
		14'h3509: color = 2'b00;
		14'h350a: color = 2'b00;
		14'h350b: color = 2'b00;
		14'h350c: color = 2'b00;
		14'h350d: color = 2'b00;
		14'h350e: color = 2'b00;
		14'h350f: color = 2'b00;
		14'h3510: color = 2'b00;
		14'h3511: color = 2'b00;
		14'h3512: color = 2'b00;
		14'h3513: color = 2'b00;
		14'h3514: color = 2'b00;
		14'h3515: color = 2'b00;
		14'h3516: color = 2'b00;
		14'h3517: color = 2'b00;
		14'h3518: color = 2'b00;
		14'h3519: color = 2'b00;
		14'h351a: color = 2'b00;
		14'h351b: color = 2'b00;
		14'h351c: color = 2'b00;
		14'h351d: color = 2'b00;
		14'h351e: color = 2'b00;
		14'h351f: color = 2'b00;
		14'h3520: color = 2'b00;
		14'h3521: color = 2'b00;
		14'h3522: color = 2'b00;
		14'h3523: color = 2'b00;
		14'h3524: color = 2'b00;
		14'h3525: color = 2'b00;
		14'h3526: color = 2'b00;
		14'h3527: color = 2'b00;
		14'h3528: color = 2'b00;
		14'h3529: color = 2'b00;
		14'h352a: color = 2'b00;
		14'h352b: color = 2'b00;
		14'h352c: color = 2'b00;
		14'h352d: color = 2'b00;
		14'h352e: color = 2'b00;
		14'h352f: color = 2'b00;
		14'h3530: color = 2'b00;
		14'h3531: color = 2'b00;
		14'h3532: color = 2'b00;
		14'h3533: color = 2'b00;
		14'h3534: color = 2'b01;
		14'h3535: color = 2'b10;
		14'h3536: color = 2'b10;
		14'h3537: color = 2'b11;
		14'h3538: color = 2'b11;
		14'h3539: color = 2'b11;
		14'h353a: color = 2'b11;
		14'h353b: color = 2'b11;
		14'h353c: color = 2'b11;
		14'h353d: color = 2'b11;
		14'h353e: color = 2'b11;
		14'h353f: color = 2'b11;
		14'h3540: color = 2'b11;
		14'h3541: color = 2'b11;
		14'h3542: color = 2'b11;
		14'h3543: color = 2'b10;
		14'h3544: color = 2'b10;
		14'h3545: color = 2'b10;
		14'h3546: color = 2'b10;
		14'h3547: color = 2'b01;
		14'h3548: color = 2'b01;
		14'h3549: color = 2'b01;
		14'h354a: color = 2'b01;
		14'h354b: color = 2'b10;
		14'h354c: color = 2'b11;
		14'h354d: color = 2'b11;
		14'h354e: color = 2'b11;
		14'h354f: color = 2'b10;
		14'h3550: color = 2'b11;
		14'h3551: color = 2'b11;
		14'h3552: color = 2'b00;
		14'h3553: color = 2'b00;
		14'h3554: color = 2'b00;
		14'h3555: color = 2'b00;
		14'h3556: color = 2'b00;
		14'h3557: color = 2'b00;
		14'h3558: color = 2'b00;
		14'h3559: color = 2'b00;
		14'h355a: color = 2'b00;
		14'h355b: color = 2'b00;
		14'h355c: color = 2'b00;
		14'h355d: color = 2'b00;
		14'h355e: color = 2'b00;
		14'h355f: color = 2'b00;
		14'h3560: color = 2'b00;
		14'h3561: color = 2'b00;
		14'h3562: color = 2'b00;
		14'h3563: color = 2'b00;
		14'h3564: color = 2'b00;
		14'h3565: color = 2'b00;
		14'h3566: color = 2'b00;
		14'h3567: color = 2'b00;
		14'h3568: color = 2'b00;
		14'h3569: color = 2'b00;
		14'h356a: color = 2'b00;
		14'h356b: color = 2'b00;
		14'h356c: color = 2'b00;
		14'h356d: color = 2'b00;
		14'h356e: color = 2'b00;
		14'h356f: color = 2'b00;
		14'h3570: color = 2'b00;
		14'h3571: color = 2'b00;
		14'h3572: color = 2'b00;
		14'h3573: color = 2'b00;
		14'h3574: color = 2'b00;
		14'h3575: color = 2'b00;
		14'h3576: color = 2'b00;
		14'h3577: color = 2'b11;
		14'h3578: color = 2'b11;
		14'h3579: color = 2'b11;
		14'h357a: color = 2'b11;
		14'h357b: color = 2'b11;
		14'h357c: color = 2'b11;
		14'h357d: color = 2'b11;
		14'h357e: color = 2'b11;
		14'h357f: color = 2'b11;
		14'h3580: color = 2'b00;
		14'h3581: color = 2'b00;
		14'h3582: color = 2'b00;
		14'h3583: color = 2'b00;
		14'h3584: color = 2'b01;
		14'h3585: color = 2'b00;
		14'h3586: color = 2'b00;
		14'h3587: color = 2'b00;
		14'h3588: color = 2'b00;
		14'h3589: color = 2'b00;
		14'h358a: color = 2'b01;
		14'h358b: color = 2'b00;
		14'h358c: color = 2'b00;
		14'h358d: color = 2'b00;
		14'h358e: color = 2'b00;
		14'h358f: color = 2'b00;
		14'h3590: color = 2'b00;
		14'h3591: color = 2'b00;
		14'h3592: color = 2'b00;
		14'h3593: color = 2'b00;
		14'h3594: color = 2'b00;
		14'h3595: color = 2'b00;
		14'h3596: color = 2'b00;
		14'h3597: color = 2'b00;
		14'h3598: color = 2'b00;
		14'h3599: color = 2'b00;
		14'h359a: color = 2'b00;
		14'h359b: color = 2'b00;
		14'h359c: color = 2'b00;
		14'h359d: color = 2'b00;
		14'h359e: color = 2'b00;
		14'h359f: color = 2'b00;
		14'h35a0: color = 2'b00;
		14'h35a1: color = 2'b00;
		14'h35a2: color = 2'b00;
		14'h35a3: color = 2'b00;
		14'h35a4: color = 2'b00;
		14'h35a5: color = 2'b00;
		14'h35a6: color = 2'b00;
		14'h35a7: color = 2'b00;
		14'h35a8: color = 2'b00;
		14'h35a9: color = 2'b00;
		14'h35aa: color = 2'b00;
		14'h35ab: color = 2'b00;
		14'h35ac: color = 2'b00;
		14'h35ad: color = 2'b00;
		14'h35ae: color = 2'b00;
		14'h35af: color = 2'b00;
		14'h35b0: color = 2'b00;
		14'h35b1: color = 2'b00;
		14'h35b2: color = 2'b00;
		14'h35b3: color = 2'b00;
		14'h35b4: color = 2'b00;
		14'h35b5: color = 2'b10;
		14'h35b6: color = 2'b10;
		14'h35b7: color = 2'b11;
		14'h35b8: color = 2'b11;
		14'h35b9: color = 2'b11;
		14'h35ba: color = 2'b11;
		14'h35bb: color = 2'b11;
		14'h35bc: color = 2'b11;
		14'h35bd: color = 2'b11;
		14'h35be: color = 2'b11;
		14'h35bf: color = 2'b11;
		14'h35c0: color = 2'b11;
		14'h35c1: color = 2'b11;
		14'h35c2: color = 2'b10;
		14'h35c3: color = 2'b01;
		14'h35c4: color = 2'b10;
		14'h35c5: color = 2'b10;
		14'h35c6: color = 2'b10;
		14'h35c7: color = 2'b01;
		14'h35c8: color = 2'b01;
		14'h35c9: color = 2'b10;
		14'h35ca: color = 2'b01;
		14'h35cb: color = 2'b00;
		14'h35cc: color = 2'b10;
		14'h35cd: color = 2'b11;
		14'h35ce: color = 2'b11;
		14'h35cf: color = 2'b11;
		14'h35d0: color = 2'b10;
		14'h35d1: color = 2'b10;
		14'h35d2: color = 2'b01;
		14'h35d3: color = 2'b00;
		14'h35d4: color = 2'b00;
		14'h35d5: color = 2'b00;
		14'h35d6: color = 2'b00;
		14'h35d7: color = 2'b00;
		14'h35d8: color = 2'b00;
		14'h35d9: color = 2'b00;
		14'h35da: color = 2'b00;
		14'h35db: color = 2'b00;
		14'h35dc: color = 2'b00;
		14'h35dd: color = 2'b00;
		14'h35de: color = 2'b00;
		14'h35df: color = 2'b00;
		14'h35e0: color = 2'b00;
		14'h35e1: color = 2'b00;
		14'h35e2: color = 2'b00;
		14'h35e3: color = 2'b00;
		14'h35e4: color = 2'b00;
		14'h35e5: color = 2'b00;
		14'h35e6: color = 2'b00;
		14'h35e7: color = 2'b00;
		14'h35e8: color = 2'b00;
		14'h35e9: color = 2'b00;
		14'h35ea: color = 2'b00;
		14'h35eb: color = 2'b00;
		14'h35ec: color = 2'b00;
		14'h35ed: color = 2'b00;
		14'h35ee: color = 2'b00;
		14'h35ef: color = 2'b00;
		14'h35f0: color = 2'b00;
		14'h35f1: color = 2'b00;
		14'h35f2: color = 2'b00;
		14'h35f3: color = 2'b00;
		14'h35f4: color = 2'b00;
		14'h35f5: color = 2'b00;
		14'h35f6: color = 2'b00;
		14'h35f7: color = 2'b11;
		14'h35f8: color = 2'b11;
		14'h35f9: color = 2'b11;
		14'h35fa: color = 2'b11;
		14'h35fb: color = 2'b11;
		14'h35fc: color = 2'b11;
		14'h35fd: color = 2'b11;
		14'h35fe: color = 2'b11;
		14'h35ff: color = 2'b11;
		14'h3600: color = 2'b00;
		14'h3601: color = 2'b01;
		14'h3602: color = 2'b00;
		14'h3603: color = 2'b00;
		14'h3604: color = 2'b00;
		14'h3605: color = 2'b00;
		14'h3606: color = 2'b00;
		14'h3607: color = 2'b00;
		14'h3608: color = 2'b00;
		14'h3609: color = 2'b00;
		14'h360a: color = 2'b00;
		14'h360b: color = 2'b00;
		14'h360c: color = 2'b01;
		14'h360d: color = 2'b00;
		14'h360e: color = 2'b00;
		14'h360f: color = 2'b00;
		14'h3610: color = 2'b00;
		14'h3611: color = 2'b00;
		14'h3612: color = 2'b00;
		14'h3613: color = 2'b00;
		14'h3614: color = 2'b00;
		14'h3615: color = 2'b00;
		14'h3616: color = 2'b00;
		14'h3617: color = 2'b00;
		14'h3618: color = 2'b00;
		14'h3619: color = 2'b00;
		14'h361a: color = 2'b00;
		14'h361b: color = 2'b00;
		14'h361c: color = 2'b00;
		14'h361d: color = 2'b00;
		14'h361e: color = 2'b00;
		14'h361f: color = 2'b00;
		14'h3620: color = 2'b00;
		14'h3621: color = 2'b00;
		14'h3622: color = 2'b00;
		14'h3623: color = 2'b00;
		14'h3624: color = 2'b00;
		14'h3625: color = 2'b00;
		14'h3626: color = 2'b00;
		14'h3627: color = 2'b00;
		14'h3628: color = 2'b00;
		14'h3629: color = 2'b00;
		14'h362a: color = 2'b00;
		14'h362b: color = 2'b00;
		14'h362c: color = 2'b00;
		14'h362d: color = 2'b00;
		14'h362e: color = 2'b01;
		14'h362f: color = 2'b00;
		14'h3630: color = 2'b00;
		14'h3631: color = 2'b00;
		14'h3632: color = 2'b00;
		14'h3633: color = 2'b00;
		14'h3634: color = 2'b00;
		14'h3635: color = 2'b01;
		14'h3636: color = 2'b10;
		14'h3637: color = 2'b10;
		14'h3638: color = 2'b10;
		14'h3639: color = 2'b11;
		14'h363a: color = 2'b11;
		14'h363b: color = 2'b11;
		14'h363c: color = 2'b11;
		14'h363d: color = 2'b11;
		14'h363e: color = 2'b11;
		14'h363f: color = 2'b11;
		14'h3640: color = 2'b11;
		14'h3641: color = 2'b11;
		14'h3642: color = 2'b01;
		14'h3643: color = 2'b10;
		14'h3644: color = 2'b10;
		14'h3645: color = 2'b10;
		14'h3646: color = 2'b10;
		14'h3647: color = 2'b10;
		14'h3648: color = 2'b10;
		14'h3649: color = 2'b10;
		14'h364a: color = 2'b01;
		14'h364b: color = 2'b01;
		14'h364c: color = 2'b01;
		14'h364d: color = 2'b10;
		14'h364e: color = 2'b10;
		14'h364f: color = 2'b11;
		14'h3650: color = 2'b11;
		14'h3651: color = 2'b11;
		14'h3652: color = 2'b01;
		14'h3653: color = 2'b00;
		14'h3654: color = 2'b00;
		14'h3655: color = 2'b00;
		14'h3656: color = 2'b00;
		14'h3657: color = 2'b00;
		14'h3658: color = 2'b00;
		14'h3659: color = 2'b00;
		14'h365a: color = 2'b00;
		14'h365b: color = 2'b00;
		14'h365c: color = 2'b00;
		14'h365d: color = 2'b00;
		14'h365e: color = 2'b00;
		14'h365f: color = 2'b00;
		14'h3660: color = 2'b00;
		14'h3661: color = 2'b00;
		14'h3662: color = 2'b00;
		14'h3663: color = 2'b00;
		14'h3664: color = 2'b00;
		14'h3665: color = 2'b00;
		14'h3666: color = 2'b00;
		14'h3667: color = 2'b00;
		14'h3668: color = 2'b00;
		14'h3669: color = 2'b00;
		14'h366a: color = 2'b00;
		14'h366b: color = 2'b00;
		14'h366c: color = 2'b00;
		14'h366d: color = 2'b00;
		14'h366e: color = 2'b00;
		14'h366f: color = 2'b00;
		14'h3670: color = 2'b00;
		14'h3671: color = 2'b00;
		14'h3672: color = 2'b00;
		14'h3673: color = 2'b00;
		14'h3674: color = 2'b00;
		14'h3675: color = 2'b00;
		14'h3676: color = 2'b00;
		14'h3677: color = 2'b01;
		14'h3678: color = 2'b01;
		14'h3679: color = 2'b11;
		14'h367a: color = 2'b11;
		14'h367b: color = 2'b11;
		14'h367c: color = 2'b11;
		14'h367d: color = 2'b11;
		14'h367e: color = 2'b11;
		14'h367f: color = 2'b11;
		14'h3680: color = 2'b00;
		14'h3681: color = 2'b00;
		14'h3682: color = 2'b01;
		14'h3683: color = 2'b00;
		14'h3684: color = 2'b00;
		14'h3685: color = 2'b00;
		14'h3686: color = 2'b00;
		14'h3687: color = 2'b00;
		14'h3688: color = 2'b00;
		14'h3689: color = 2'b00;
		14'h368a: color = 2'b01;
		14'h368b: color = 2'b00;
		14'h368c: color = 2'b00;
		14'h368d: color = 2'b00;
		14'h368e: color = 2'b00;
		14'h368f: color = 2'b00;
		14'h3690: color = 2'b00;
		14'h3691: color = 2'b00;
		14'h3692: color = 2'b00;
		14'h3693: color = 2'b00;
		14'h3694: color = 2'b00;
		14'h3695: color = 2'b00;
		14'h3696: color = 2'b00;
		14'h3697: color = 2'b00;
		14'h3698: color = 2'b00;
		14'h3699: color = 2'b00;
		14'h369a: color = 2'b00;
		14'h369b: color = 2'b00;
		14'h369c: color = 2'b00;
		14'h369d: color = 2'b00;
		14'h369e: color = 2'b00;
		14'h369f: color = 2'b00;
		14'h36a0: color = 2'b00;
		14'h36a1: color = 2'b00;
		14'h36a2: color = 2'b00;
		14'h36a3: color = 2'b00;
		14'h36a4: color = 2'b00;
		14'h36a5: color = 2'b00;
		14'h36a6: color = 2'b00;
		14'h36a7: color = 2'b00;
		14'h36a8: color = 2'b00;
		14'h36a9: color = 2'b00;
		14'h36aa: color = 2'b00;
		14'h36ab: color = 2'b00;
		14'h36ac: color = 2'b00;
		14'h36ad: color = 2'b00;
		14'h36ae: color = 2'b00;
		14'h36af: color = 2'b00;
		14'h36b0: color = 2'b00;
		14'h36b1: color = 2'b00;
		14'h36b2: color = 2'b00;
		14'h36b3: color = 2'b00;
		14'h36b4: color = 2'b00;
		14'h36b5: color = 2'b01;
		14'h36b6: color = 2'b10;
		14'h36b7: color = 2'b10;
		14'h36b8: color = 2'b10;
		14'h36b9: color = 2'b11;
		14'h36ba: color = 2'b11;
		14'h36bb: color = 2'b11;
		14'h36bc: color = 2'b11;
		14'h36bd: color = 2'b11;
		14'h36be: color = 2'b11;
		14'h36bf: color = 2'b11;
		14'h36c0: color = 2'b10;
		14'h36c1: color = 2'b10;
		14'h36c2: color = 2'b10;
		14'h36c3: color = 2'b10;
		14'h36c4: color = 2'b10;
		14'h36c5: color = 2'b01;
		14'h36c6: color = 2'b10;
		14'h36c7: color = 2'b01;
		14'h36c8: color = 2'b01;
		14'h36c9: color = 2'b01;
		14'h36ca: color = 2'b01;
		14'h36cb: color = 2'b10;
		14'h36cc: color = 2'b01;
		14'h36cd: color = 2'b01;
		14'h36ce: color = 2'b10;
		14'h36cf: color = 2'b11;
		14'h36d0: color = 2'b10;
		14'h36d1: color = 2'b11;
		14'h36d2: color = 2'b00;
		14'h36d3: color = 2'b00;
		14'h36d4: color = 2'b00;
		14'h36d5: color = 2'b00;
		14'h36d6: color = 2'b00;
		14'h36d7: color = 2'b00;
		14'h36d8: color = 2'b00;
		14'h36d9: color = 2'b00;
		14'h36da: color = 2'b00;
		14'h36db: color = 2'b00;
		14'h36dc: color = 2'b00;
		14'h36dd: color = 2'b00;
		14'h36de: color = 2'b00;
		14'h36df: color = 2'b00;
		14'h36e0: color = 2'b00;
		14'h36e1: color = 2'b00;
		14'h36e2: color = 2'b00;
		14'h36e3: color = 2'b00;
		14'h36e4: color = 2'b00;
		14'h36e5: color = 2'b00;
		14'h36e6: color = 2'b00;
		14'h36e7: color = 2'b00;
		14'h36e8: color = 2'b00;
		14'h36e9: color = 2'b00;
		14'h36ea: color = 2'b00;
		14'h36eb: color = 2'b00;
		14'h36ec: color = 2'b00;
		14'h36ed: color = 2'b00;
		14'h36ee: color = 2'b00;
		14'h36ef: color = 2'b00;
		14'h36f0: color = 2'b00;
		14'h36f1: color = 2'b00;
		14'h36f2: color = 2'b00;
		14'h36f3: color = 2'b00;
		14'h36f4: color = 2'b00;
		14'h36f5: color = 2'b00;
		14'h36f6: color = 2'b00;
		14'h36f7: color = 2'b00;
		14'h36f8: color = 2'b00;
		14'h36f9: color = 2'b11;
		14'h36fa: color = 2'b11;
		14'h36fb: color = 2'b11;
		14'h36fc: color = 2'b11;
		14'h36fd: color = 2'b11;
		14'h36fe: color = 2'b11;
		14'h36ff: color = 2'b11;
		14'h3700: color = 2'b00;
		14'h3701: color = 2'b00;
		14'h3702: color = 2'b00;
		14'h3703: color = 2'b00;
		14'h3704: color = 2'b00;
		14'h3705: color = 2'b00;
		14'h3706: color = 2'b00;
		14'h3707: color = 2'b00;
		14'h3708: color = 2'b00;
		14'h3709: color = 2'b00;
		14'h370a: color = 2'b00;
		14'h370b: color = 2'b00;
		14'h370c: color = 2'b00;
		14'h370d: color = 2'b00;
		14'h370e: color = 2'b00;
		14'h370f: color = 2'b00;
		14'h3710: color = 2'b00;
		14'h3711: color = 2'b00;
		14'h3712: color = 2'b00;
		14'h3713: color = 2'b00;
		14'h3714: color = 2'b00;
		14'h3715: color = 2'b00;
		14'h3716: color = 2'b00;
		14'h3717: color = 2'b00;
		14'h3718: color = 2'b00;
		14'h3719: color = 2'b00;
		14'h371a: color = 2'b00;
		14'h371b: color = 2'b00;
		14'h371c: color = 2'b00;
		14'h371d: color = 2'b00;
		14'h371e: color = 2'b00;
		14'h371f: color = 2'b00;
		14'h3720: color = 2'b00;
		14'h3721: color = 2'b00;
		14'h3722: color = 2'b00;
		14'h3723: color = 2'b00;
		14'h3724: color = 2'b00;
		14'h3725: color = 2'b00;
		14'h3726: color = 2'b00;
		14'h3727: color = 2'b00;
		14'h3728: color = 2'b00;
		14'h3729: color = 2'b00;
		14'h372a: color = 2'b00;
		14'h372b: color = 2'b00;
		14'h372c: color = 2'b00;
		14'h372d: color = 2'b00;
		14'h372e: color = 2'b00;
		14'h372f: color = 2'b00;
		14'h3730: color = 2'b00;
		14'h3731: color = 2'b00;
		14'h3732: color = 2'b00;
		14'h3733: color = 2'b00;
		14'h3734: color = 2'b00;
		14'h3735: color = 2'b00;
		14'h3736: color = 2'b10;
		14'h3737: color = 2'b10;
		14'h3738: color = 2'b10;
		14'h3739: color = 2'b10;
		14'h373a: color = 2'b11;
		14'h373b: color = 2'b11;
		14'h373c: color = 2'b11;
		14'h373d: color = 2'b11;
		14'h373e: color = 2'b11;
		14'h373f: color = 2'b10;
		14'h3740: color = 2'b01;
		14'h3741: color = 2'b10;
		14'h3742: color = 2'b10;
		14'h3743: color = 2'b10;
		14'h3744: color = 2'b10;
		14'h3745: color = 2'b01;
		14'h3746: color = 2'b10;
		14'h3747: color = 2'b10;
		14'h3748: color = 2'b10;
		14'h3749: color = 2'b01;
		14'h374a: color = 2'b10;
		14'h374b: color = 2'b10;
		14'h374c: color = 2'b01;
		14'h374d: color = 2'b00;
		14'h374e: color = 2'b01;
		14'h374f: color = 2'b11;
		14'h3750: color = 2'b10;
		14'h3751: color = 2'b11;
		14'h3752: color = 2'b01;
		14'h3753: color = 2'b00;
		14'h3754: color = 2'b00;
		14'h3755: color = 2'b00;
		14'h3756: color = 2'b00;
		14'h3757: color = 2'b00;
		14'h3758: color = 2'b00;
		14'h3759: color = 2'b00;
		14'h375a: color = 2'b00;
		14'h375b: color = 2'b00;
		14'h375c: color = 2'b00;
		14'h375d: color = 2'b00;
		14'h375e: color = 2'b00;
		14'h375f: color = 2'b00;
		14'h3760: color = 2'b00;
		14'h3761: color = 2'b00;
		14'h3762: color = 2'b00;
		14'h3763: color = 2'b00;
		14'h3764: color = 2'b00;
		14'h3765: color = 2'b00;
		14'h3766: color = 2'b00;
		14'h3767: color = 2'b00;
		14'h3768: color = 2'b00;
		14'h3769: color = 2'b00;
		14'h376a: color = 2'b00;
		14'h376b: color = 2'b00;
		14'h376c: color = 2'b00;
		14'h376d: color = 2'b00;
		14'h376e: color = 2'b00;
		14'h376f: color = 2'b00;
		14'h3770: color = 2'b00;
		14'h3771: color = 2'b00;
		14'h3772: color = 2'b00;
		14'h3773: color = 2'b00;
		14'h3774: color = 2'b00;
		14'h3775: color = 2'b00;
		14'h3776: color = 2'b00;
		14'h3777: color = 2'b00;
		14'h3778: color = 2'b00;
		14'h3779: color = 2'b11;
		14'h377a: color = 2'b11;
		14'h377b: color = 2'b11;
		14'h377c: color = 2'b11;
		14'h377d: color = 2'b11;
		14'h377e: color = 2'b11;
		14'h377f: color = 2'b11;
		14'h3780: color = 2'b01;
		14'h3781: color = 2'b00;
		14'h3782: color = 2'b00;
		14'h3783: color = 2'b00;
		14'h3784: color = 2'b00;
		14'h3785: color = 2'b00;
		14'h3786: color = 2'b01;
		14'h3787: color = 2'b00;
		14'h3788: color = 2'b00;
		14'h3789: color = 2'b00;
		14'h378a: color = 2'b00;
		14'h378b: color = 2'b00;
		14'h378c: color = 2'b00;
		14'h378d: color = 2'b00;
		14'h378e: color = 2'b00;
		14'h378f: color = 2'b00;
		14'h3790: color = 2'b00;
		14'h3791: color = 2'b00;
		14'h3792: color = 2'b00;
		14'h3793: color = 2'b00;
		14'h3794: color = 2'b00;
		14'h3795: color = 2'b00;
		14'h3796: color = 2'b00;
		14'h3797: color = 2'b00;
		14'h3798: color = 2'b00;
		14'h3799: color = 2'b00;
		14'h379a: color = 2'b00;
		14'h379b: color = 2'b00;
		14'h379c: color = 2'b00;
		14'h379d: color = 2'b00;
		14'h379e: color = 2'b00;
		14'h379f: color = 2'b00;
		14'h37a0: color = 2'b00;
		14'h37a1: color = 2'b00;
		14'h37a2: color = 2'b00;
		14'h37a3: color = 2'b00;
		14'h37a4: color = 2'b00;
		14'h37a5: color = 2'b00;
		14'h37a6: color = 2'b00;
		14'h37a7: color = 2'b00;
		14'h37a8: color = 2'b00;
		14'h37a9: color = 2'b00;
		14'h37aa: color = 2'b00;
		14'h37ab: color = 2'b00;
		14'h37ac: color = 2'b00;
		14'h37ad: color = 2'b00;
		14'h37ae: color = 2'b00;
		14'h37af: color = 2'b00;
		14'h37b0: color = 2'b00;
		14'h37b1: color = 2'b00;
		14'h37b2: color = 2'b00;
		14'h37b3: color = 2'b00;
		14'h37b4: color = 2'b00;
		14'h37b5: color = 2'b00;
		14'h37b6: color = 2'b01;
		14'h37b7: color = 2'b10;
		14'h37b8: color = 2'b10;
		14'h37b9: color = 2'b11;
		14'h37ba: color = 2'b10;
		14'h37bb: color = 2'b11;
		14'h37bc: color = 2'b11;
		14'h37bd: color = 2'b11;
		14'h37be: color = 2'b01;
		14'h37bf: color = 2'b00;
		14'h37c0: color = 2'b01;
		14'h37c1: color = 2'b10;
		14'h37c2: color = 2'b10;
		14'h37c3: color = 2'b10;
		14'h37c4: color = 2'b10;
		14'h37c5: color = 2'b10;
		14'h37c6: color = 2'b10;
		14'h37c7: color = 2'b10;
		14'h37c8: color = 2'b10;
		14'h37c9: color = 2'b10;
		14'h37ca: color = 2'b01;
		14'h37cb: color = 2'b10;
		14'h37cc: color = 2'b01;
		14'h37cd: color = 2'b01;
		14'h37ce: color = 2'b00;
		14'h37cf: color = 2'b10;
		14'h37d0: color = 2'b11;
		14'h37d1: color = 2'b11;
		14'h37d2: color = 2'b01;
		14'h37d3: color = 2'b00;
		14'h37d4: color = 2'b00;
		14'h37d5: color = 2'b00;
		14'h37d6: color = 2'b00;
		14'h37d7: color = 2'b00;
		14'h37d8: color = 2'b00;
		14'h37d9: color = 2'b00;
		14'h37da: color = 2'b00;
		14'h37db: color = 2'b00;
		14'h37dc: color = 2'b00;
		14'h37dd: color = 2'b00;
		14'h37de: color = 2'b00;
		14'h37df: color = 2'b00;
		14'h37e0: color = 2'b00;
		14'h37e1: color = 2'b00;
		14'h37e2: color = 2'b00;
		14'h37e3: color = 2'b00;
		14'h37e4: color = 2'b00;
		14'h37e5: color = 2'b00;
		14'h37e6: color = 2'b00;
		14'h37e7: color = 2'b00;
		14'h37e8: color = 2'b00;
		14'h37e9: color = 2'b00;
		14'h37ea: color = 2'b00;
		14'h37eb: color = 2'b00;
		14'h37ec: color = 2'b00;
		14'h37ed: color = 2'b00;
		14'h37ee: color = 2'b00;
		14'h37ef: color = 2'b00;
		14'h37f0: color = 2'b00;
		14'h37f1: color = 2'b00;
		14'h37f2: color = 2'b00;
		14'h37f3: color = 2'b00;
		14'h37f4: color = 2'b00;
		14'h37f5: color = 2'b00;
		14'h37f6: color = 2'b00;
		14'h37f7: color = 2'b00;
		14'h37f8: color = 2'b00;
		14'h37f9: color = 2'b11;
		14'h37fa: color = 2'b11;
		14'h37fb: color = 2'b11;
		14'h37fc: color = 2'b11;
		14'h37fd: color = 2'b11;
		14'h37fe: color = 2'b11;
		14'h37ff: color = 2'b11;
		14'h3800: color = 2'b00;
		14'h3801: color = 2'b00;
		14'h3802: color = 2'b00;
		14'h3803: color = 2'b01;
		14'h3804: color = 2'b00;
		14'h3805: color = 2'b00;
		14'h3806: color = 2'b01;
		14'h3807: color = 2'b00;
		14'h3808: color = 2'b00;
		14'h3809: color = 2'b00;
		14'h380a: color = 2'b00;
		14'h380b: color = 2'b00;
		14'h380c: color = 2'b00;
		14'h380d: color = 2'b00;
		14'h380e: color = 2'b00;
		14'h380f: color = 2'b00;
		14'h3810: color = 2'b00;
		14'h3811: color = 2'b00;
		14'h3812: color = 2'b00;
		14'h3813: color = 2'b00;
		14'h3814: color = 2'b00;
		14'h3815: color = 2'b00;
		14'h3816: color = 2'b00;
		14'h3817: color = 2'b00;
		14'h3818: color = 2'b00;
		14'h3819: color = 2'b00;
		14'h381a: color = 2'b00;
		14'h381b: color = 2'b00;
		14'h381c: color = 2'b00;
		14'h381d: color = 2'b00;
		14'h381e: color = 2'b00;
		14'h381f: color = 2'b00;
		14'h3820: color = 2'b00;
		14'h3821: color = 2'b00;
		14'h3822: color = 2'b00;
		14'h3823: color = 2'b00;
		14'h3824: color = 2'b00;
		14'h3825: color = 2'b00;
		14'h3826: color = 2'b00;
		14'h3827: color = 2'b00;
		14'h3828: color = 2'b00;
		14'h3829: color = 2'b00;
		14'h382a: color = 2'b00;
		14'h382b: color = 2'b00;
		14'h382c: color = 2'b00;
		14'h382d: color = 2'b00;
		14'h382e: color = 2'b00;
		14'h382f: color = 2'b00;
		14'h3830: color = 2'b00;
		14'h3831: color = 2'b00;
		14'h3832: color = 2'b00;
		14'h3833: color = 2'b00;
		14'h3834: color = 2'b00;
		14'h3835: color = 2'b00;
		14'h3836: color = 2'b00;
		14'h3837: color = 2'b10;
		14'h3838: color = 2'b10;
		14'h3839: color = 2'b11;
		14'h383a: color = 2'b10;
		14'h383b: color = 2'b11;
		14'h383c: color = 2'b11;
		14'h383d: color = 2'b10;
		14'h383e: color = 2'b00;
		14'h383f: color = 2'b00;
		14'h3840: color = 2'b00;
		14'h3841: color = 2'b10;
		14'h3842: color = 2'b10;
		14'h3843: color = 2'b11;
		14'h3844: color = 2'b10;
		14'h3845: color = 2'b10;
		14'h3846: color = 2'b10;
		14'h3847: color = 2'b10;
		14'h3848: color = 2'b10;
		14'h3849: color = 2'b10;
		14'h384a: color = 2'b10;
		14'h384b: color = 2'b10;
		14'h384c: color = 2'b01;
		14'h384d: color = 2'b01;
		14'h384e: color = 2'b00;
		14'h384f: color = 2'b01;
		14'h3850: color = 2'b11;
		14'h3851: color = 2'b11;
		14'h3852: color = 2'b01;
		14'h3853: color = 2'b00;
		14'h3854: color = 2'b00;
		14'h3855: color = 2'b00;
		14'h3856: color = 2'b00;
		14'h3857: color = 2'b00;
		14'h3858: color = 2'b00;
		14'h3859: color = 2'b00;
		14'h385a: color = 2'b00;
		14'h385b: color = 2'b00;
		14'h385c: color = 2'b00;
		14'h385d: color = 2'b00;
		14'h385e: color = 2'b00;
		14'h385f: color = 2'b00;
		14'h3860: color = 2'b00;
		14'h3861: color = 2'b00;
		14'h3862: color = 2'b00;
		14'h3863: color = 2'b00;
		14'h3864: color = 2'b00;
		14'h3865: color = 2'b00;
		14'h3866: color = 2'b00;
		14'h3867: color = 2'b00;
		14'h3868: color = 2'b00;
		14'h3869: color = 2'b00;
		14'h386a: color = 2'b00;
		14'h386b: color = 2'b00;
		14'h386c: color = 2'b00;
		14'h386d: color = 2'b00;
		14'h386e: color = 2'b00;
		14'h386f: color = 2'b00;
		14'h3870: color = 2'b00;
		14'h3871: color = 2'b00;
		14'h3872: color = 2'b00;
		14'h3873: color = 2'b00;
		14'h3874: color = 2'b00;
		14'h3875: color = 2'b00;
		14'h3876: color = 2'b00;
		14'h3877: color = 2'b00;
		14'h3878: color = 2'b00;
		14'h3879: color = 2'b01;
		14'h387a: color = 2'b11;
		14'h387b: color = 2'b11;
		14'h387c: color = 2'b11;
		14'h387d: color = 2'b11;
		14'h387e: color = 2'b11;
		14'h387f: color = 2'b11;
		14'h3880: color = 2'b00;
		14'h3881: color = 2'b00;
		14'h3882: color = 2'b00;
		14'h3883: color = 2'b00;
		14'h3884: color = 2'b00;
		14'h3885: color = 2'b00;
		14'h3886: color = 2'b00;
		14'h3887: color = 2'b00;
		14'h3888: color = 2'b00;
		14'h3889: color = 2'b01;
		14'h388a: color = 2'b00;
		14'h388b: color = 2'b00;
		14'h388c: color = 2'b00;
		14'h388d: color = 2'b00;
		14'h388e: color = 2'b00;
		14'h388f: color = 2'b00;
		14'h3890: color = 2'b00;
		14'h3891: color = 2'b00;
		14'h3892: color = 2'b00;
		14'h3893: color = 2'b00;
		14'h3894: color = 2'b00;
		14'h3895: color = 2'b00;
		14'h3896: color = 2'b00;
		14'h3897: color = 2'b00;
		14'h3898: color = 2'b00;
		14'h3899: color = 2'b00;
		14'h389a: color = 2'b00;
		14'h389b: color = 2'b00;
		14'h389c: color = 2'b00;
		14'h389d: color = 2'b00;
		14'h389e: color = 2'b00;
		14'h389f: color = 2'b00;
		14'h38a0: color = 2'b00;
		14'h38a1: color = 2'b00;
		14'h38a2: color = 2'b00;
		14'h38a3: color = 2'b00;
		14'h38a4: color = 2'b00;
		14'h38a5: color = 2'b00;
		14'h38a6: color = 2'b00;
		14'h38a7: color = 2'b00;
		14'h38a8: color = 2'b00;
		14'h38a9: color = 2'b00;
		14'h38aa: color = 2'b00;
		14'h38ab: color = 2'b00;
		14'h38ac: color = 2'b00;
		14'h38ad: color = 2'b00;
		14'h38ae: color = 2'b00;
		14'h38af: color = 2'b00;
		14'h38b0: color = 2'b00;
		14'h38b1: color = 2'b00;
		14'h38b2: color = 2'b00;
		14'h38b3: color = 2'b00;
		14'h38b4: color = 2'b00;
		14'h38b5: color = 2'b00;
		14'h38b6: color = 2'b00;
		14'h38b7: color = 2'b01;
		14'h38b8: color = 2'b01;
		14'h38b9: color = 2'b10;
		14'h38ba: color = 2'b11;
		14'h38bb: color = 2'b10;
		14'h38bc: color = 2'b10;
		14'h38bd: color = 2'b10;
		14'h38be: color = 2'b00;
		14'h38bf: color = 2'b01;
		14'h38c0: color = 2'b00;
		14'h38c1: color = 2'b01;
		14'h38c2: color = 2'b10;
		14'h38c3: color = 2'b10;
		14'h38c4: color = 2'b11;
		14'h38c5: color = 2'b10;
		14'h38c6: color = 2'b11;
		14'h38c7: color = 2'b10;
		14'h38c8: color = 2'b10;
		14'h38c9: color = 2'b10;
		14'h38ca: color = 2'b10;
		14'h38cb: color = 2'b10;
		14'h38cc: color = 2'b01;
		14'h38cd: color = 2'b01;
		14'h38ce: color = 2'b01;
		14'h38cf: color = 2'b01;
		14'h38d0: color = 2'b10;
		14'h38d1: color = 2'b11;
		14'h38d2: color = 2'b01;
		14'h38d3: color = 2'b00;
		14'h38d4: color = 2'b00;
		14'h38d5: color = 2'b00;
		14'h38d6: color = 2'b00;
		14'h38d7: color = 2'b00;
		14'h38d8: color = 2'b00;
		14'h38d9: color = 2'b00;
		14'h38da: color = 2'b00;
		14'h38db: color = 2'b00;
		14'h38dc: color = 2'b00;
		14'h38dd: color = 2'b00;
		14'h38de: color = 2'b00;
		14'h38df: color = 2'b00;
		14'h38e0: color = 2'b00;
		14'h38e1: color = 2'b00;
		14'h38e2: color = 2'b00;
		14'h38e3: color = 2'b00;
		14'h38e4: color = 2'b00;
		14'h38e5: color = 2'b00;
		14'h38e6: color = 2'b00;
		14'h38e7: color = 2'b00;
		14'h38e8: color = 2'b00;
		14'h38e9: color = 2'b00;
		14'h38ea: color = 2'b00;
		14'h38eb: color = 2'b00;
		14'h38ec: color = 2'b00;
		14'h38ed: color = 2'b00;
		14'h38ee: color = 2'b00;
		14'h38ef: color = 2'b00;
		14'h38f0: color = 2'b00;
		14'h38f1: color = 2'b00;
		14'h38f2: color = 2'b00;
		14'h38f3: color = 2'b00;
		14'h38f4: color = 2'b00;
		14'h38f5: color = 2'b00;
		14'h38f6: color = 2'b00;
		14'h38f7: color = 2'b00;
		14'h38f8: color = 2'b00;
		14'h38f9: color = 2'b00;
		14'h38fa: color = 2'b11;
		14'h38fb: color = 2'b11;
		14'h38fc: color = 2'b11;
		14'h38fd: color = 2'b11;
		14'h38fe: color = 2'b11;
		14'h38ff: color = 2'b11;
		14'h3900: color = 2'b00;
		14'h3901: color = 2'b00;
		14'h3902: color = 2'b00;
		14'h3903: color = 2'b01;
		14'h3904: color = 2'b00;
		14'h3905: color = 2'b00;
		14'h3906: color = 2'b00;
		14'h3907: color = 2'b00;
		14'h3908: color = 2'b00;
		14'h3909: color = 2'b00;
		14'h390a: color = 2'b00;
		14'h390b: color = 2'b00;
		14'h390c: color = 2'b00;
		14'h390d: color = 2'b00;
		14'h390e: color = 2'b00;
		14'h390f: color = 2'b00;
		14'h3910: color = 2'b00;
		14'h3911: color = 2'b00;
		14'h3912: color = 2'b00;
		14'h3913: color = 2'b00;
		14'h3914: color = 2'b00;
		14'h3915: color = 2'b00;
		14'h3916: color = 2'b00;
		14'h3917: color = 2'b00;
		14'h3918: color = 2'b00;
		14'h3919: color = 2'b00;
		14'h391a: color = 2'b00;
		14'h391b: color = 2'b00;
		14'h391c: color = 2'b00;
		14'h391d: color = 2'b00;
		14'h391e: color = 2'b00;
		14'h391f: color = 2'b00;
		14'h3920: color = 2'b00;
		14'h3921: color = 2'b00;
		14'h3922: color = 2'b00;
		14'h3923: color = 2'b00;
		14'h3924: color = 2'b00;
		14'h3925: color = 2'b00;
		14'h3926: color = 2'b00;
		14'h3927: color = 2'b00;
		14'h3928: color = 2'b00;
		14'h3929: color = 2'b00;
		14'h392a: color = 2'b00;
		14'h392b: color = 2'b00;
		14'h392c: color = 2'b00;
		14'h392d: color = 2'b00;
		14'h392e: color = 2'b00;
		14'h392f: color = 2'b00;
		14'h3930: color = 2'b00;
		14'h3931: color = 2'b00;
		14'h3932: color = 2'b00;
		14'h3933: color = 2'b00;
		14'h3934: color = 2'b00;
		14'h3935: color = 2'b00;
		14'h3936: color = 2'b00;
		14'h3937: color = 2'b00;
		14'h3938: color = 2'b00;
		14'h3939: color = 2'b11;
		14'h393a: color = 2'b10;
		14'h393b: color = 2'b10;
		14'h393c: color = 2'b10;
		14'h393d: color = 2'b11;
		14'h393e: color = 2'b01;
		14'h393f: color = 2'b00;
		14'h3940: color = 2'b00;
		14'h3941: color = 2'b00;
		14'h3942: color = 2'b01;
		14'h3943: color = 2'b11;
		14'h3944: color = 2'b11;
		14'h3945: color = 2'b10;
		14'h3946: color = 2'b10;
		14'h3947: color = 2'b10;
		14'h3948: color = 2'b10;
		14'h3949: color = 2'b10;
		14'h394a: color = 2'b11;
		14'h394b: color = 2'b10;
		14'h394c: color = 2'b01;
		14'h394d: color = 2'b10;
		14'h394e: color = 2'b10;
		14'h394f: color = 2'b10;
		14'h3950: color = 2'b10;
		14'h3951: color = 2'b11;
		14'h3952: color = 2'b01;
		14'h3953: color = 2'b00;
		14'h3954: color = 2'b00;
		14'h3955: color = 2'b00;
		14'h3956: color = 2'b00;
		14'h3957: color = 2'b00;
		14'h3958: color = 2'b00;
		14'h3959: color = 2'b00;
		14'h395a: color = 2'b00;
		14'h395b: color = 2'b00;
		14'h395c: color = 2'b00;
		14'h395d: color = 2'b00;
		14'h395e: color = 2'b00;
		14'h395f: color = 2'b00;
		14'h3960: color = 2'b00;
		14'h3961: color = 2'b00;
		14'h3962: color = 2'b00;
		14'h3963: color = 2'b00;
		14'h3964: color = 2'b00;
		14'h3965: color = 2'b00;
		14'h3966: color = 2'b00;
		14'h3967: color = 2'b00;
		14'h3968: color = 2'b00;
		14'h3969: color = 2'b00;
		14'h396a: color = 2'b00;
		14'h396b: color = 2'b00;
		14'h396c: color = 2'b00;
		14'h396d: color = 2'b00;
		14'h396e: color = 2'b00;
		14'h396f: color = 2'b00;
		14'h3970: color = 2'b00;
		14'h3971: color = 2'b00;
		14'h3972: color = 2'b00;
		14'h3973: color = 2'b00;
		14'h3974: color = 2'b00;
		14'h3975: color = 2'b00;
		14'h3976: color = 2'b00;
		14'h3977: color = 2'b00;
		14'h3978: color = 2'b00;
		14'h3979: color = 2'b00;
		14'h397a: color = 2'b11;
		14'h397b: color = 2'b11;
		14'h397c: color = 2'b11;
		14'h397d: color = 2'b11;
		14'h397e: color = 2'b11;
		14'h397f: color = 2'b11;
		14'h3980: color = 2'b00;
		14'h3981: color = 2'b00;
		14'h3982: color = 2'b00;
		14'h3983: color = 2'b00;
		14'h3984: color = 2'b01;
		14'h3985: color = 2'b00;
		14'h3986: color = 2'b00;
		14'h3987: color = 2'b00;
		14'h3988: color = 2'b00;
		14'h3989: color = 2'b00;
		14'h398a: color = 2'b00;
		14'h398b: color = 2'b00;
		14'h398c: color = 2'b00;
		14'h398d: color = 2'b00;
		14'h398e: color = 2'b00;
		14'h398f: color = 2'b00;
		14'h3990: color = 2'b00;
		14'h3991: color = 2'b00;
		14'h3992: color = 2'b00;
		14'h3993: color = 2'b00;
		14'h3994: color = 2'b00;
		14'h3995: color = 2'b00;
		14'h3996: color = 2'b00;
		14'h3997: color = 2'b00;
		14'h3998: color = 2'b00;
		14'h3999: color = 2'b00;
		14'h399a: color = 2'b00;
		14'h399b: color = 2'b00;
		14'h399c: color = 2'b00;
		14'h399d: color = 2'b00;
		14'h399e: color = 2'b00;
		14'h399f: color = 2'b00;
		14'h39a0: color = 2'b00;
		14'h39a1: color = 2'b00;
		14'h39a2: color = 2'b00;
		14'h39a3: color = 2'b00;
		14'h39a4: color = 2'b00;
		14'h39a5: color = 2'b00;
		14'h39a6: color = 2'b00;
		14'h39a7: color = 2'b00;
		14'h39a8: color = 2'b00;
		14'h39a9: color = 2'b00;
		14'h39aa: color = 2'b00;
		14'h39ab: color = 2'b00;
		14'h39ac: color = 2'b00;
		14'h39ad: color = 2'b00;
		14'h39ae: color = 2'b00;
		14'h39af: color = 2'b00;
		14'h39b0: color = 2'b00;
		14'h39b1: color = 2'b00;
		14'h39b2: color = 2'b00;
		14'h39b3: color = 2'b00;
		14'h39b4: color = 2'b00;
		14'h39b5: color = 2'b00;
		14'h39b6: color = 2'b00;
		14'h39b7: color = 2'b00;
		14'h39b8: color = 2'b00;
		14'h39b9: color = 2'b01;
		14'h39ba: color = 2'b10;
		14'h39bb: color = 2'b10;
		14'h39bc: color = 2'b10;
		14'h39bd: color = 2'b11;
		14'h39be: color = 2'b10;
		14'h39bf: color = 2'b00;
		14'h39c0: color = 2'b01;
		14'h39c1: color = 2'b01;
		14'h39c2: color = 2'b00;
		14'h39c3: color = 2'b10;
		14'h39c4: color = 2'b10;
		14'h39c5: color = 2'b10;
		14'h39c6: color = 2'b10;
		14'h39c7: color = 2'b11;
		14'h39c8: color = 2'b11;
		14'h39c9: color = 2'b10;
		14'h39ca: color = 2'b10;
		14'h39cb: color = 2'b10;
		14'h39cc: color = 2'b01;
		14'h39cd: color = 2'b10;
		14'h39ce: color = 2'b11;
		14'h39cf: color = 2'b10;
		14'h39d0: color = 2'b10;
		14'h39d1: color = 2'b11;
		14'h39d2: color = 2'b10;
		14'h39d3: color = 2'b00;
		14'h39d4: color = 2'b00;
		14'h39d5: color = 2'b00;
		14'h39d6: color = 2'b00;
		14'h39d7: color = 2'b00;
		14'h39d8: color = 2'b00;
		14'h39d9: color = 2'b00;
		14'h39da: color = 2'b00;
		14'h39db: color = 2'b00;
		14'h39dc: color = 2'b00;
		14'h39dd: color = 2'b00;
		14'h39de: color = 2'b00;
		14'h39df: color = 2'b00;
		14'h39e0: color = 2'b00;
		14'h39e1: color = 2'b00;
		14'h39e2: color = 2'b00;
		14'h39e3: color = 2'b00;
		14'h39e4: color = 2'b00;
		14'h39e5: color = 2'b00;
		14'h39e6: color = 2'b00;
		14'h39e7: color = 2'b00;
		14'h39e8: color = 2'b00;
		14'h39e9: color = 2'b00;
		14'h39ea: color = 2'b00;
		14'h39eb: color = 2'b00;
		14'h39ec: color = 2'b00;
		14'h39ed: color = 2'b00;
		14'h39ee: color = 2'b00;
		14'h39ef: color = 2'b00;
		14'h39f0: color = 2'b00;
		14'h39f1: color = 2'b00;
		14'h39f2: color = 2'b00;
		14'h39f3: color = 2'b00;
		14'h39f4: color = 2'b00;
		14'h39f5: color = 2'b00;
		14'h39f6: color = 2'b00;
		14'h39f7: color = 2'b00;
		14'h39f8: color = 2'b00;
		14'h39f9: color = 2'b00;
		14'h39fa: color = 2'b11;
		14'h39fb: color = 2'b11;
		14'h39fc: color = 2'b11;
		14'h39fd: color = 2'b11;
		14'h39fe: color = 2'b11;
		14'h39ff: color = 2'b11;
		14'h3a00: color = 2'b00;
		14'h3a01: color = 2'b00;
		14'h3a02: color = 2'b00;
		14'h3a03: color = 2'b00;
		14'h3a04: color = 2'b00;
		14'h3a05: color = 2'b00;
		14'h3a06: color = 2'b00;
		14'h3a07: color = 2'b00;
		14'h3a08: color = 2'b00;
		14'h3a09: color = 2'b00;
		14'h3a0a: color = 2'b00;
		14'h3a0b: color = 2'b00;
		14'h3a0c: color = 2'b00;
		14'h3a0d: color = 2'b00;
		14'h3a0e: color = 2'b00;
		14'h3a0f: color = 2'b00;
		14'h3a10: color = 2'b00;
		14'h3a11: color = 2'b00;
		14'h3a12: color = 2'b00;
		14'h3a13: color = 2'b00;
		14'h3a14: color = 2'b00;
		14'h3a15: color = 2'b00;
		14'h3a16: color = 2'b00;
		14'h3a17: color = 2'b00;
		14'h3a18: color = 2'b00;
		14'h3a19: color = 2'b00;
		14'h3a1a: color = 2'b00;
		14'h3a1b: color = 2'b00;
		14'h3a1c: color = 2'b00;
		14'h3a1d: color = 2'b00;
		14'h3a1e: color = 2'b00;
		14'h3a1f: color = 2'b00;
		14'h3a20: color = 2'b00;
		14'h3a21: color = 2'b00;
		14'h3a22: color = 2'b00;
		14'h3a23: color = 2'b00;
		14'h3a24: color = 2'b00;
		14'h3a25: color = 2'b00;
		14'h3a26: color = 2'b00;
		14'h3a27: color = 2'b00;
		14'h3a28: color = 2'b00;
		14'h3a29: color = 2'b00;
		14'h3a2a: color = 2'b00;
		14'h3a2b: color = 2'b00;
		14'h3a2c: color = 2'b00;
		14'h3a2d: color = 2'b00;
		14'h3a2e: color = 2'b00;
		14'h3a2f: color = 2'b00;
		14'h3a30: color = 2'b00;
		14'h3a31: color = 2'b00;
		14'h3a32: color = 2'b00;
		14'h3a33: color = 2'b00;
		14'h3a34: color = 2'b00;
		14'h3a35: color = 2'b00;
		14'h3a36: color = 2'b00;
		14'h3a37: color = 2'b00;
		14'h3a38: color = 2'b00;
		14'h3a39: color = 2'b01;
		14'h3a3a: color = 2'b11;
		14'h3a3b: color = 2'b11;
		14'h3a3c: color = 2'b10;
		14'h3a3d: color = 2'b11;
		14'h3a3e: color = 2'b11;
		14'h3a3f: color = 2'b01;
		14'h3a40: color = 2'b01;
		14'h3a41: color = 2'b01;
		14'h3a42: color = 2'b00;
		14'h3a43: color = 2'b01;
		14'h3a44: color = 2'b10;
		14'h3a45: color = 2'b10;
		14'h3a46: color = 2'b11;
		14'h3a47: color = 2'b10;
		14'h3a48: color = 2'b10;
		14'h3a49: color = 2'b11;
		14'h3a4a: color = 2'b11;
		14'h3a4b: color = 2'b10;
		14'h3a4c: color = 2'b10;
		14'h3a4d: color = 2'b10;
		14'h3a4e: color = 2'b10;
		14'h3a4f: color = 2'b11;
		14'h3a50: color = 2'b10;
		14'h3a51: color = 2'b10;
		14'h3a52: color = 2'b10;
		14'h3a53: color = 2'b00;
		14'h3a54: color = 2'b00;
		14'h3a55: color = 2'b00;
		14'h3a56: color = 2'b00;
		14'h3a57: color = 2'b00;
		14'h3a58: color = 2'b00;
		14'h3a59: color = 2'b00;
		14'h3a5a: color = 2'b00;
		14'h3a5b: color = 2'b00;
		14'h3a5c: color = 2'b00;
		14'h3a5d: color = 2'b00;
		14'h3a5e: color = 2'b00;
		14'h3a5f: color = 2'b00;
		14'h3a60: color = 2'b00;
		14'h3a61: color = 2'b00;
		14'h3a62: color = 2'b00;
		14'h3a63: color = 2'b00;
		14'h3a64: color = 2'b00;
		14'h3a65: color = 2'b00;
		14'h3a66: color = 2'b00;
		14'h3a67: color = 2'b00;
		14'h3a68: color = 2'b00;
		14'h3a69: color = 2'b00;
		14'h3a6a: color = 2'b00;
		14'h3a6b: color = 2'b00;
		14'h3a6c: color = 2'b00;
		14'h3a6d: color = 2'b00;
		14'h3a6e: color = 2'b00;
		14'h3a6f: color = 2'b00;
		14'h3a70: color = 2'b00;
		14'h3a71: color = 2'b00;
		14'h3a72: color = 2'b00;
		14'h3a73: color = 2'b00;
		14'h3a74: color = 2'b00;
		14'h3a75: color = 2'b00;
		14'h3a76: color = 2'b00;
		14'h3a77: color = 2'b00;
		14'h3a78: color = 2'b00;
		14'h3a79: color = 2'b00;
		14'h3a7a: color = 2'b11;
		14'h3a7b: color = 2'b11;
		14'h3a7c: color = 2'b11;
		14'h3a7d: color = 2'b11;
		14'h3a7e: color = 2'b11;
		14'h3a7f: color = 2'b11;
		14'h3a80: color = 2'b00;
		14'h3a81: color = 2'b00;
		14'h3a82: color = 2'b00;
		14'h3a83: color = 2'b00;
		14'h3a84: color = 2'b00;
		14'h3a85: color = 2'b00;
		14'h3a86: color = 2'b00;
		14'h3a87: color = 2'b00;
		14'h3a88: color = 2'b00;
		14'h3a89: color = 2'b00;
		14'h3a8a: color = 2'b00;
		14'h3a8b: color = 2'b00;
		14'h3a8c: color = 2'b00;
		14'h3a8d: color = 2'b00;
		14'h3a8e: color = 2'b00;
		14'h3a8f: color = 2'b00;
		14'h3a90: color = 2'b00;
		14'h3a91: color = 2'b00;
		14'h3a92: color = 2'b00;
		14'h3a93: color = 2'b00;
		14'h3a94: color = 2'b00;
		14'h3a95: color = 2'b00;
		14'h3a96: color = 2'b00;
		14'h3a97: color = 2'b00;
		14'h3a98: color = 2'b00;
		14'h3a99: color = 2'b00;
		14'h3a9a: color = 2'b00;
		14'h3a9b: color = 2'b00;
		14'h3a9c: color = 2'b00;
		14'h3a9d: color = 2'b00;
		14'h3a9e: color = 2'b00;
		14'h3a9f: color = 2'b00;
		14'h3aa0: color = 2'b00;
		14'h3aa1: color = 2'b00;
		14'h3aa2: color = 2'b00;
		14'h3aa3: color = 2'b00;
		14'h3aa4: color = 2'b00;
		14'h3aa5: color = 2'b00;
		14'h3aa6: color = 2'b00;
		14'h3aa7: color = 2'b00;
		14'h3aa8: color = 2'b00;
		14'h3aa9: color = 2'b00;
		14'h3aaa: color = 2'b00;
		14'h3aab: color = 2'b00;
		14'h3aac: color = 2'b00;
		14'h3aad: color = 2'b00;
		14'h3aae: color = 2'b00;
		14'h3aaf: color = 2'b01;
		14'h3ab0: color = 2'b00;
		14'h3ab1: color = 2'b00;
		14'h3ab2: color = 2'b00;
		14'h3ab3: color = 2'b00;
		14'h3ab4: color = 2'b00;
		14'h3ab5: color = 2'b00;
		14'h3ab6: color = 2'b00;
		14'h3ab7: color = 2'b00;
		14'h3ab8: color = 2'b00;
		14'h3ab9: color = 2'b00;
		14'h3aba: color = 2'b10;
		14'h3abb: color = 2'b11;
		14'h3abc: color = 2'b11;
		14'h3abd: color = 2'b10;
		14'h3abe: color = 2'b11;
		14'h3abf: color = 2'b11;
		14'h3ac0: color = 2'b10;
		14'h3ac1: color = 2'b01;
		14'h3ac2: color = 2'b01;
		14'h3ac3: color = 2'b00;
		14'h3ac4: color = 2'b01;
		14'h3ac5: color = 2'b10;
		14'h3ac6: color = 2'b10;
		14'h3ac7: color = 2'b10;
		14'h3ac8: color = 2'b10;
		14'h3ac9: color = 2'b10;
		14'h3aca: color = 2'b10;
		14'h3acb: color = 2'b11;
		14'h3acc: color = 2'b01;
		14'h3acd: color = 2'b10;
		14'h3ace: color = 2'b11;
		14'h3acf: color = 2'b11;
		14'h3ad0: color = 2'b11;
		14'h3ad1: color = 2'b10;
		14'h3ad2: color = 2'b10;
		14'h3ad3: color = 2'b00;
		14'h3ad4: color = 2'b00;
		14'h3ad5: color = 2'b00;
		14'h3ad6: color = 2'b00;
		14'h3ad7: color = 2'b00;
		14'h3ad8: color = 2'b00;
		14'h3ad9: color = 2'b00;
		14'h3ada: color = 2'b00;
		14'h3adb: color = 2'b00;
		14'h3adc: color = 2'b00;
		14'h3add: color = 2'b00;
		14'h3ade: color = 2'b00;
		14'h3adf: color = 2'b00;
		14'h3ae0: color = 2'b00;
		14'h3ae1: color = 2'b00;
		14'h3ae2: color = 2'b00;
		14'h3ae3: color = 2'b00;
		14'h3ae4: color = 2'b00;
		14'h3ae5: color = 2'b00;
		14'h3ae6: color = 2'b00;
		14'h3ae7: color = 2'b00;
		14'h3ae8: color = 2'b00;
		14'h3ae9: color = 2'b00;
		14'h3aea: color = 2'b00;
		14'h3aeb: color = 2'b00;
		14'h3aec: color = 2'b00;
		14'h3aed: color = 2'b00;
		14'h3aee: color = 2'b00;
		14'h3aef: color = 2'b00;
		14'h3af0: color = 2'b00;
		14'h3af1: color = 2'b00;
		14'h3af2: color = 2'b00;
		14'h3af3: color = 2'b00;
		14'h3af4: color = 2'b00;
		14'h3af5: color = 2'b00;
		14'h3af6: color = 2'b00;
		14'h3af7: color = 2'b00;
		14'h3af8: color = 2'b00;
		14'h3af9: color = 2'b00;
		14'h3afa: color = 2'b11;
		14'h3afb: color = 2'b11;
		14'h3afc: color = 2'b11;
		14'h3afd: color = 2'b11;
		14'h3afe: color = 2'b11;
		14'h3aff: color = 2'b11;
		14'h3b00: color = 2'b00;
		14'h3b01: color = 2'b01;
		14'h3b02: color = 2'b00;
		14'h3b03: color = 2'b00;
		14'h3b04: color = 2'b00;
		14'h3b05: color = 2'b00;
		14'h3b06: color = 2'b00;
		14'h3b07: color = 2'b00;
		14'h3b08: color = 2'b00;
		14'h3b09: color = 2'b00;
		14'h3b0a: color = 2'b00;
		14'h3b0b: color = 2'b00;
		14'h3b0c: color = 2'b00;
		14'h3b0d: color = 2'b00;
		14'h3b0e: color = 2'b00;
		14'h3b0f: color = 2'b00;
		14'h3b10: color = 2'b00;
		14'h3b11: color = 2'b00;
		14'h3b12: color = 2'b00;
		14'h3b13: color = 2'b00;
		14'h3b14: color = 2'b00;
		14'h3b15: color = 2'b00;
		14'h3b16: color = 2'b00;
		14'h3b17: color = 2'b00;
		14'h3b18: color = 2'b00;
		14'h3b19: color = 2'b00;
		14'h3b1a: color = 2'b00;
		14'h3b1b: color = 2'b00;
		14'h3b1c: color = 2'b00;
		14'h3b1d: color = 2'b00;
		14'h3b1e: color = 2'b00;
		14'h3b1f: color = 2'b00;
		14'h3b20: color = 2'b00;
		14'h3b21: color = 2'b00;
		14'h3b22: color = 2'b00;
		14'h3b23: color = 2'b00;
		14'h3b24: color = 2'b00;
		14'h3b25: color = 2'b00;
		14'h3b26: color = 2'b00;
		14'h3b27: color = 2'b00;
		14'h3b28: color = 2'b00;
		14'h3b29: color = 2'b00;
		14'h3b2a: color = 2'b00;
		14'h3b2b: color = 2'b00;
		14'h3b2c: color = 2'b00;
		14'h3b2d: color = 2'b00;
		14'h3b2e: color = 2'b00;
		14'h3b2f: color = 2'b00;
		14'h3b30: color = 2'b00;
		14'h3b31: color = 2'b00;
		14'h3b32: color = 2'b00;
		14'h3b33: color = 2'b00;
		14'h3b34: color = 2'b00;
		14'h3b35: color = 2'b00;
		14'h3b36: color = 2'b00;
		14'h3b37: color = 2'b00;
		14'h3b38: color = 2'b00;
		14'h3b39: color = 2'b00;
		14'h3b3a: color = 2'b01;
		14'h3b3b: color = 2'b11;
		14'h3b3c: color = 2'b11;
		14'h3b3d: color = 2'b11;
		14'h3b3e: color = 2'b11;
		14'h3b3f: color = 2'b10;
		14'h3b40: color = 2'b10;
		14'h3b41: color = 2'b10;
		14'h3b42: color = 2'b01;
		14'h3b43: color = 2'b01;
		14'h3b44: color = 2'b01;
		14'h3b45: color = 2'b01;
		14'h3b46: color = 2'b10;
		14'h3b47: color = 2'b11;
		14'h3b48: color = 2'b11;
		14'h3b49: color = 2'b10;
		14'h3b4a: color = 2'b10;
		14'h3b4b: color = 2'b10;
		14'h3b4c: color = 2'b10;
		14'h3b4d: color = 2'b10;
		14'h3b4e: color = 2'b11;
		14'h3b4f: color = 2'b11;
		14'h3b50: color = 2'b10;
		14'h3b51: color = 2'b11;
		14'h3b52: color = 2'b10;
		14'h3b53: color = 2'b01;
		14'h3b54: color = 2'b00;
		14'h3b55: color = 2'b00;
		14'h3b56: color = 2'b00;
		14'h3b57: color = 2'b00;
		14'h3b58: color = 2'b00;
		14'h3b59: color = 2'b00;
		14'h3b5a: color = 2'b00;
		14'h3b5b: color = 2'b00;
		14'h3b5c: color = 2'b00;
		14'h3b5d: color = 2'b00;
		14'h3b5e: color = 2'b00;
		14'h3b5f: color = 2'b00;
		14'h3b60: color = 2'b00;
		14'h3b61: color = 2'b00;
		14'h3b62: color = 2'b00;
		14'h3b63: color = 2'b00;
		14'h3b64: color = 2'b00;
		14'h3b65: color = 2'b00;
		14'h3b66: color = 2'b00;
		14'h3b67: color = 2'b00;
		14'h3b68: color = 2'b00;
		14'h3b69: color = 2'b00;
		14'h3b6a: color = 2'b00;
		14'h3b6b: color = 2'b00;
		14'h3b6c: color = 2'b00;
		14'h3b6d: color = 2'b00;
		14'h3b6e: color = 2'b00;
		14'h3b6f: color = 2'b00;
		14'h3b70: color = 2'b00;
		14'h3b71: color = 2'b00;
		14'h3b72: color = 2'b00;
		14'h3b73: color = 2'b00;
		14'h3b74: color = 2'b00;
		14'h3b75: color = 2'b00;
		14'h3b76: color = 2'b00;
		14'h3b77: color = 2'b00;
		14'h3b78: color = 2'b00;
		14'h3b79: color = 2'b00;
		14'h3b7a: color = 2'b11;
		14'h3b7b: color = 2'b11;
		14'h3b7c: color = 2'b11;
		14'h3b7d: color = 2'b11;
		14'h3b7e: color = 2'b11;
		14'h3b7f: color = 2'b11;
		14'h3b80: color = 2'b00;
		14'h3b81: color = 2'b00;
		14'h3b82: color = 2'b00;
		14'h3b83: color = 2'b00;
		14'h3b84: color = 2'b00;
		14'h3b85: color = 2'b00;
		14'h3b86: color = 2'b00;
		14'h3b87: color = 2'b00;
		14'h3b88: color = 2'b00;
		14'h3b89: color = 2'b00;
		14'h3b8a: color = 2'b00;
		14'h3b8b: color = 2'b00;
		14'h3b8c: color = 2'b00;
		14'h3b8d: color = 2'b00;
		14'h3b8e: color = 2'b00;
		14'h3b8f: color = 2'b00;
		14'h3b90: color = 2'b00;
		14'h3b91: color = 2'b00;
		14'h3b92: color = 2'b00;
		14'h3b93: color = 2'b00;
		14'h3b94: color = 2'b00;
		14'h3b95: color = 2'b00;
		14'h3b96: color = 2'b00;
		14'h3b97: color = 2'b00;
		14'h3b98: color = 2'b00;
		14'h3b99: color = 2'b00;
		14'h3b9a: color = 2'b00;
		14'h3b9b: color = 2'b00;
		14'h3b9c: color = 2'b00;
		14'h3b9d: color = 2'b00;
		14'h3b9e: color = 2'b00;
		14'h3b9f: color = 2'b00;
		14'h3ba0: color = 2'b00;
		14'h3ba1: color = 2'b00;
		14'h3ba2: color = 2'b00;
		14'h3ba3: color = 2'b00;
		14'h3ba4: color = 2'b00;
		14'h3ba5: color = 2'b00;
		14'h3ba6: color = 2'b00;
		14'h3ba7: color = 2'b00;
		14'h3ba8: color = 2'b00;
		14'h3ba9: color = 2'b00;
		14'h3baa: color = 2'b00;
		14'h3bab: color = 2'b00;
		14'h3bac: color = 2'b00;
		14'h3bad: color = 2'b00;
		14'h3bae: color = 2'b00;
		14'h3baf: color = 2'b00;
		14'h3bb0: color = 2'b00;
		14'h3bb1: color = 2'b00;
		14'h3bb2: color = 2'b00;
		14'h3bb3: color = 2'b00;
		14'h3bb4: color = 2'b00;
		14'h3bb5: color = 2'b00;
		14'h3bb6: color = 2'b00;
		14'h3bb7: color = 2'b00;
		14'h3bb8: color = 2'b00;
		14'h3bb9: color = 2'b00;
		14'h3bba: color = 2'b00;
		14'h3bbb: color = 2'b10;
		14'h3bbc: color = 2'b11;
		14'h3bbd: color = 2'b11;
		14'h3bbe: color = 2'b11;
		14'h3bbf: color = 2'b11;
		14'h3bc0: color = 2'b11;
		14'h3bc1: color = 2'b11;
		14'h3bc2: color = 2'b10;
		14'h3bc3: color = 2'b01;
		14'h3bc4: color = 2'b00;
		14'h3bc5: color = 2'b01;
		14'h3bc6: color = 2'b10;
		14'h3bc7: color = 2'b11;
		14'h3bc8: color = 2'b11;
		14'h3bc9: color = 2'b10;
		14'h3bca: color = 2'b11;
		14'h3bcb: color = 2'b10;
		14'h3bcc: color = 2'b10;
		14'h3bcd: color = 2'b10;
		14'h3bce: color = 2'b10;
		14'h3bcf: color = 2'b11;
		14'h3bd0: color = 2'b11;
		14'h3bd1: color = 2'b11;
		14'h3bd2: color = 2'b10;
		14'h3bd3: color = 2'b01;
		14'h3bd4: color = 2'b00;
		14'h3bd5: color = 2'b00;
		14'h3bd6: color = 2'b00;
		14'h3bd7: color = 2'b00;
		14'h3bd8: color = 2'b00;
		14'h3bd9: color = 2'b00;
		14'h3bda: color = 2'b00;
		14'h3bdb: color = 2'b00;
		14'h3bdc: color = 2'b00;
		14'h3bdd: color = 2'b00;
		14'h3bde: color = 2'b00;
		14'h3bdf: color = 2'b00;
		14'h3be0: color = 2'b00;
		14'h3be1: color = 2'b00;
		14'h3be2: color = 2'b00;
		14'h3be3: color = 2'b00;
		14'h3be4: color = 2'b00;
		14'h3be5: color = 2'b00;
		14'h3be6: color = 2'b00;
		14'h3be7: color = 2'b00;
		14'h3be8: color = 2'b00;
		14'h3be9: color = 2'b00;
		14'h3bea: color = 2'b00;
		14'h3beb: color = 2'b00;
		14'h3bec: color = 2'b00;
		14'h3bed: color = 2'b00;
		14'h3bee: color = 2'b00;
		14'h3bef: color = 2'b00;
		14'h3bf0: color = 2'b00;
		14'h3bf1: color = 2'b00;
		14'h3bf2: color = 2'b00;
		14'h3bf3: color = 2'b00;
		14'h3bf4: color = 2'b00;
		14'h3bf5: color = 2'b00;
		14'h3bf6: color = 2'b00;
		14'h3bf7: color = 2'b00;
		14'h3bf8: color = 2'b00;
		14'h3bf9: color = 2'b00;
		14'h3bfa: color = 2'b11;
		14'h3bfb: color = 2'b11;
		14'h3bfc: color = 2'b11;
		14'h3bfd: color = 2'b11;
		14'h3bfe: color = 2'b11;
		14'h3bff: color = 2'b11;
		14'h3c00: color = 2'b00;
		14'h3c01: color = 2'b00;
		14'h3c02: color = 2'b00;
		14'h3c03: color = 2'b00;
		14'h3c04: color = 2'b00;
		14'h3c05: color = 2'b00;
		14'h3c06: color = 2'b00;
		14'h3c07: color = 2'b00;
		14'h3c08: color = 2'b00;
		14'h3c09: color = 2'b00;
		14'h3c0a: color = 2'b00;
		14'h3c0b: color = 2'b00;
		14'h3c0c: color = 2'b00;
		14'h3c0d: color = 2'b00;
		14'h3c0e: color = 2'b00;
		14'h3c0f: color = 2'b00;
		14'h3c10: color = 2'b00;
		14'h3c11: color = 2'b00;
		14'h3c12: color = 2'b00;
		14'h3c13: color = 2'b00;
		14'h3c14: color = 2'b00;
		14'h3c15: color = 2'b00;
		14'h3c16: color = 2'b00;
		14'h3c17: color = 2'b00;
		14'h3c18: color = 2'b00;
		14'h3c19: color = 2'b00;
		14'h3c1a: color = 2'b00;
		14'h3c1b: color = 2'b00;
		14'h3c1c: color = 2'b00;
		14'h3c1d: color = 2'b00;
		14'h3c1e: color = 2'b00;
		14'h3c1f: color = 2'b00;
		14'h3c20: color = 2'b00;
		14'h3c21: color = 2'b00;
		14'h3c22: color = 2'b00;
		14'h3c23: color = 2'b00;
		14'h3c24: color = 2'b00;
		14'h3c25: color = 2'b00;
		14'h3c26: color = 2'b00;
		14'h3c27: color = 2'b00;
		14'h3c28: color = 2'b00;
		14'h3c29: color = 2'b00;
		14'h3c2a: color = 2'b00;
		14'h3c2b: color = 2'b00;
		14'h3c2c: color = 2'b00;
		14'h3c2d: color = 2'b00;
		14'h3c2e: color = 2'b00;
		14'h3c2f: color = 2'b00;
		14'h3c30: color = 2'b00;
		14'h3c31: color = 2'b00;
		14'h3c32: color = 2'b00;
		14'h3c33: color = 2'b00;
		14'h3c34: color = 2'b00;
		14'h3c35: color = 2'b00;
		14'h3c36: color = 2'b00;
		14'h3c37: color = 2'b00;
		14'h3c38: color = 2'b00;
		14'h3c39: color = 2'b00;
		14'h3c3a: color = 2'b00;
		14'h3c3b: color = 2'b10;
		14'h3c3c: color = 2'b11;
		14'h3c3d: color = 2'b11;
		14'h3c3e: color = 2'b11;
		14'h3c3f: color = 2'b11;
		14'h3c40: color = 2'b11;
		14'h3c41: color = 2'b11;
		14'h3c42: color = 2'b10;
		14'h3c43: color = 2'b01;
		14'h3c44: color = 2'b00;
		14'h3c45: color = 2'b01;
		14'h3c46: color = 2'b10;
		14'h3c47: color = 2'b11;
		14'h3c48: color = 2'b11;
		14'h3c49: color = 2'b10;
		14'h3c4a: color = 2'b11;
		14'h3c4b: color = 2'b10;
		14'h3c4c: color = 2'b10;
		14'h3c4d: color = 2'b10;
		14'h3c4e: color = 2'b10;
		14'h3c4f: color = 2'b11;
		14'h3c50: color = 2'b11;
		14'h3c51: color = 2'b11;
		14'h3c52: color = 2'b10;
		14'h3c53: color = 2'b01;
		14'h3c54: color = 2'b00;
		14'h3c55: color = 2'b00;
		14'h3c56: color = 2'b00;
		14'h3c57: color = 2'b00;
		14'h3c58: color = 2'b00;
		14'h3c59: color = 2'b00;
		14'h3c5a: color = 2'b00;
		14'h3c5b: color = 2'b00;
		14'h3c5c: color = 2'b00;
		14'h3c5d: color = 2'b00;
		14'h3c5e: color = 2'b00;
		14'h3c5f: color = 2'b00;
		14'h3c60: color = 2'b00;
		14'h3c61: color = 2'b00;
		14'h3c62: color = 2'b00;
		14'h3c63: color = 2'b00;
		14'h3c64: color = 2'b00;
		14'h3c65: color = 2'b00;
		14'h3c66: color = 2'b00;
		14'h3c67: color = 2'b00;
		14'h3c68: color = 2'b00;
		14'h3c69: color = 2'b00;
		14'h3c6a: color = 2'b00;
		14'h3c6b: color = 2'b00;
		14'h3c6c: color = 2'b00;
		14'h3c6d: color = 2'b00;
		14'h3c6e: color = 2'b00;
		14'h3c6f: color = 2'b00;
		14'h3c70: color = 2'b00;
		14'h3c71: color = 2'b00;
		14'h3c72: color = 2'b00;
		14'h3c73: color = 2'b00;
		14'h3c74: color = 2'b00;
		14'h3c75: color = 2'b00;
		14'h3c76: color = 2'b00;
		14'h3c77: color = 2'b00;
		14'h3c78: color = 2'b00;
		14'h3c79: color = 2'b00;
		14'h3c7a: color = 2'b11;
		14'h3c7b: color = 2'b11;
		14'h3c7c: color = 2'b11;
		14'h3c7d: color = 2'b11;
		14'h3c7e: color = 2'b11;
		14'h3c7f: color = 2'b11;
		14'h3c80: color = 2'b00;
		14'h3c81: color = 2'b00;
		14'h3c82: color = 2'b00;
		14'h3c83: color = 2'b00;
		14'h3c84: color = 2'b00;
		14'h3c85: color = 2'b00;
		14'h3c86: color = 2'b00;
		14'h3c87: color = 2'b00;
		14'h3c88: color = 2'b00;
		14'h3c89: color = 2'b00;
		14'h3c8a: color = 2'b00;
		14'h3c8b: color = 2'b00;
		14'h3c8c: color = 2'b00;
		14'h3c8d: color = 2'b00;
		14'h3c8e: color = 2'b00;
		14'h3c8f: color = 2'b00;
		14'h3c90: color = 2'b00;
		14'h3c91: color = 2'b00;
		14'h3c92: color = 2'b00;
		14'h3c93: color = 2'b00;
		14'h3c94: color = 2'b00;
		14'h3c95: color = 2'b00;
		14'h3c96: color = 2'b00;
		14'h3c97: color = 2'b00;
		14'h3c98: color = 2'b00;
		14'h3c99: color = 2'b00;
		14'h3c9a: color = 2'b00;
		14'h3c9b: color = 2'b00;
		14'h3c9c: color = 2'b00;
		14'h3c9d: color = 2'b00;
		14'h3c9e: color = 2'b00;
		14'h3c9f: color = 2'b00;
		14'h3ca0: color = 2'b00;
		14'h3ca1: color = 2'b00;
		14'h3ca2: color = 2'b00;
		14'h3ca3: color = 2'b00;
		14'h3ca4: color = 2'b00;
		14'h3ca5: color = 2'b00;
		14'h3ca6: color = 2'b00;
		14'h3ca7: color = 2'b00;
		14'h3ca8: color = 2'b00;
		14'h3ca9: color = 2'b00;
		14'h3caa: color = 2'b00;
		14'h3cab: color = 2'b00;
		14'h3cac: color = 2'b00;
		14'h3cad: color = 2'b00;
		14'h3cae: color = 2'b00;
		14'h3caf: color = 2'b00;
		14'h3cb0: color = 2'b00;
		14'h3cb1: color = 2'b00;
		14'h3cb2: color = 2'b00;
		14'h3cb3: color = 2'b00;
		14'h3cb4: color = 2'b00;
		14'h3cb5: color = 2'b00;
		14'h3cb6: color = 2'b00;
		14'h3cb7: color = 2'b00;
		14'h3cb8: color = 2'b00;
		14'h3cb9: color = 2'b00;
		14'h3cba: color = 2'b00;
		14'h3cbb: color = 2'b01;
		14'h3cbc: color = 2'b11;
		14'h3cbd: color = 2'b11;
		14'h3cbe: color = 2'b11;
		14'h3cbf: color = 2'b11;
		14'h3cc0: color = 2'b11;
		14'h3cc1: color = 2'b11;
		14'h3cc2: color = 2'b10;
		14'h3cc3: color = 2'b01;
		14'h3cc4: color = 2'b01;
		14'h3cc5: color = 2'b01;
		14'h3cc6: color = 2'b10;
		14'h3cc7: color = 2'b10;
		14'h3cc8: color = 2'b10;
		14'h3cc9: color = 2'b11;
		14'h3cca: color = 2'b10;
		14'h3ccb: color = 2'b10;
		14'h3ccc: color = 2'b10;
		14'h3ccd: color = 2'b10;
		14'h3cce: color = 2'b11;
		14'h3ccf: color = 2'b11;
		14'h3cd0: color = 2'b11;
		14'h3cd1: color = 2'b11;
		14'h3cd2: color = 2'b11;
		14'h3cd3: color = 2'b01;
		14'h3cd4: color = 2'b00;
		14'h3cd5: color = 2'b00;
		14'h3cd6: color = 2'b00;
		14'h3cd7: color = 2'b00;
		14'h3cd8: color = 2'b00;
		14'h3cd9: color = 2'b00;
		14'h3cda: color = 2'b00;
		14'h3cdb: color = 2'b00;
		14'h3cdc: color = 2'b00;
		14'h3cdd: color = 2'b00;
		14'h3cde: color = 2'b00;
		14'h3cdf: color = 2'b00;
		14'h3ce0: color = 2'b00;
		14'h3ce1: color = 2'b00;
		14'h3ce2: color = 2'b00;
		14'h3ce3: color = 2'b00;
		14'h3ce4: color = 2'b00;
		14'h3ce5: color = 2'b00;
		14'h3ce6: color = 2'b00;
		14'h3ce7: color = 2'b00;
		14'h3ce8: color = 2'b00;
		14'h3ce9: color = 2'b00;
		14'h3cea: color = 2'b00;
		14'h3ceb: color = 2'b00;
		14'h3cec: color = 2'b00;
		14'h3ced: color = 2'b00;
		14'h3cee: color = 2'b00;
		14'h3cef: color = 2'b00;
		14'h3cf0: color = 2'b00;
		14'h3cf1: color = 2'b00;
		14'h3cf2: color = 2'b00;
		14'h3cf3: color = 2'b00;
		14'h3cf4: color = 2'b00;
		14'h3cf5: color = 2'b00;
		14'h3cf6: color = 2'b00;
		14'h3cf7: color = 2'b00;
		14'h3cf8: color = 2'b00;
		14'h3cf9: color = 2'b00;
		14'h3cfa: color = 2'b10;
		14'h3cfb: color = 2'b11;
		14'h3cfc: color = 2'b11;
		14'h3cfd: color = 2'b11;
		14'h3cfe: color = 2'b11;
		14'h3cff: color = 2'b11;
		14'h3d00: color = 2'b00;
		14'h3d01: color = 2'b01;
		14'h3d02: color = 2'b00;
		14'h3d03: color = 2'b00;
		14'h3d04: color = 2'b00;
		14'h3d05: color = 2'b00;
		14'h3d06: color = 2'b00;
		14'h3d07: color = 2'b00;
		14'h3d08: color = 2'b00;
		14'h3d09: color = 2'b00;
		14'h3d0a: color = 2'b00;
		14'h3d0b: color = 2'b00;
		14'h3d0c: color = 2'b00;
		14'h3d0d: color = 2'b00;
		14'h3d0e: color = 2'b00;
		14'h3d0f: color = 2'b00;
		14'h3d10: color = 2'b00;
		14'h3d11: color = 2'b00;
		14'h3d12: color = 2'b00;
		14'h3d13: color = 2'b00;
		14'h3d14: color = 2'b00;
		14'h3d15: color = 2'b00;
		14'h3d16: color = 2'b00;
		14'h3d17: color = 2'b00;
		14'h3d18: color = 2'b00;
		14'h3d19: color = 2'b00;
		14'h3d1a: color = 2'b00;
		14'h3d1b: color = 2'b00;
		14'h3d1c: color = 2'b00;
		14'h3d1d: color = 2'b00;
		14'h3d1e: color = 2'b00;
		14'h3d1f: color = 2'b00;
		14'h3d20: color = 2'b00;
		14'h3d21: color = 2'b00;
		14'h3d22: color = 2'b00;
		14'h3d23: color = 2'b00;
		14'h3d24: color = 2'b00;
		14'h3d25: color = 2'b00;
		14'h3d26: color = 2'b00;
		14'h3d27: color = 2'b00;
		14'h3d28: color = 2'b00;
		14'h3d29: color = 2'b00;
		14'h3d2a: color = 2'b00;
		14'h3d2b: color = 2'b00;
		14'h3d2c: color = 2'b00;
		14'h3d2d: color = 2'b00;
		14'h3d2e: color = 2'b00;
		14'h3d2f: color = 2'b00;
		14'h3d30: color = 2'b00;
		14'h3d31: color = 2'b00;
		14'h3d32: color = 2'b00;
		14'h3d33: color = 2'b00;
		14'h3d34: color = 2'b00;
		14'h3d35: color = 2'b00;
		14'h3d36: color = 2'b00;
		14'h3d37: color = 2'b00;
		14'h3d38: color = 2'b00;
		14'h3d39: color = 2'b00;
		14'h3d3a: color = 2'b00;
		14'h3d3b: color = 2'b00;
		14'h3d3c: color = 2'b10;
		14'h3d3d: color = 2'b11;
		14'h3d3e: color = 2'b11;
		14'h3d3f: color = 2'b10;
		14'h3d40: color = 2'b11;
		14'h3d41: color = 2'b11;
		14'h3d42: color = 2'b11;
		14'h3d43: color = 2'b01;
		14'h3d44: color = 2'b01;
		14'h3d45: color = 2'b00;
		14'h3d46: color = 2'b10;
		14'h3d47: color = 2'b10;
		14'h3d48: color = 2'b10;
		14'h3d49: color = 2'b11;
		14'h3d4a: color = 2'b10;
		14'h3d4b: color = 2'b10;
		14'h3d4c: color = 2'b01;
		14'h3d4d: color = 2'b10;
		14'h3d4e: color = 2'b11;
		14'h3d4f: color = 2'b11;
		14'h3d50: color = 2'b11;
		14'h3d51: color = 2'b10;
		14'h3d52: color = 2'b11;
		14'h3d53: color = 2'b01;
		14'h3d54: color = 2'b01;
		14'h3d55: color = 2'b00;
		14'h3d56: color = 2'b00;
		14'h3d57: color = 2'b00;
		14'h3d58: color = 2'b00;
		14'h3d59: color = 2'b00;
		14'h3d5a: color = 2'b00;
		14'h3d5b: color = 2'b00;
		14'h3d5c: color = 2'b00;
		14'h3d5d: color = 2'b00;
		14'h3d5e: color = 2'b00;
		14'h3d5f: color = 2'b00;
		14'h3d60: color = 2'b00;
		14'h3d61: color = 2'b00;
		14'h3d62: color = 2'b00;
		14'h3d63: color = 2'b00;
		14'h3d64: color = 2'b00;
		14'h3d65: color = 2'b00;
		14'h3d66: color = 2'b00;
		14'h3d67: color = 2'b00;
		14'h3d68: color = 2'b00;
		14'h3d69: color = 2'b00;
		14'h3d6a: color = 2'b00;
		14'h3d6b: color = 2'b00;
		14'h3d6c: color = 2'b00;
		14'h3d6d: color = 2'b00;
		14'h3d6e: color = 2'b00;
		14'h3d6f: color = 2'b00;
		14'h3d70: color = 2'b00;
		14'h3d71: color = 2'b00;
		14'h3d72: color = 2'b00;
		14'h3d73: color = 2'b00;
		14'h3d74: color = 2'b00;
		14'h3d75: color = 2'b00;
		14'h3d76: color = 2'b00;
		14'h3d77: color = 2'b00;
		14'h3d78: color = 2'b00;
		14'h3d79: color = 2'b00;
		14'h3d7a: color = 2'b01;
		14'h3d7b: color = 2'b11;
		14'h3d7c: color = 2'b11;
		14'h3d7d: color = 2'b11;
		14'h3d7e: color = 2'b11;
		14'h3d7f: color = 2'b11;
		14'h3d80: color = 2'b00;
		14'h3d81: color = 2'b00;
		14'h3d82: color = 2'b01;
		14'h3d83: color = 2'b00;
		14'h3d84: color = 2'b00;
		14'h3d85: color = 2'b00;
		14'h3d86: color = 2'b00;
		14'h3d87: color = 2'b00;
		14'h3d88: color = 2'b00;
		14'h3d89: color = 2'b00;
		14'h3d8a: color = 2'b00;
		14'h3d8b: color = 2'b00;
		14'h3d8c: color = 2'b00;
		14'h3d8d: color = 2'b00;
		14'h3d8e: color = 2'b00;
		14'h3d8f: color = 2'b00;
		14'h3d90: color = 2'b00;
		14'h3d91: color = 2'b00;
		14'h3d92: color = 2'b00;
		14'h3d93: color = 2'b00;
		14'h3d94: color = 2'b00;
		14'h3d95: color = 2'b00;
		14'h3d96: color = 2'b00;
		14'h3d97: color = 2'b00;
		14'h3d98: color = 2'b00;
		14'h3d99: color = 2'b00;
		14'h3d9a: color = 2'b00;
		14'h3d9b: color = 2'b00;
		14'h3d9c: color = 2'b00;
		14'h3d9d: color = 2'b00;
		14'h3d9e: color = 2'b00;
		14'h3d9f: color = 2'b00;
		14'h3da0: color = 2'b00;
		14'h3da1: color = 2'b00;
		14'h3da2: color = 2'b00;
		14'h3da3: color = 2'b00;
		14'h3da4: color = 2'b00;
		14'h3da5: color = 2'b00;
		14'h3da6: color = 2'b00;
		14'h3da7: color = 2'b00;
		14'h3da8: color = 2'b00;
		14'h3da9: color = 2'b00;
		14'h3daa: color = 2'b00;
		14'h3dab: color = 2'b00;
		14'h3dac: color = 2'b00;
		14'h3dad: color = 2'b00;
		14'h3dae: color = 2'b00;
		14'h3daf: color = 2'b00;
		14'h3db0: color = 2'b00;
		14'h3db1: color = 2'b00;
		14'h3db2: color = 2'b00;
		14'h3db3: color = 2'b00;
		14'h3db4: color = 2'b00;
		14'h3db5: color = 2'b00;
		14'h3db6: color = 2'b00;
		14'h3db7: color = 2'b00;
		14'h3db8: color = 2'b00;
		14'h3db9: color = 2'b00;
		14'h3dba: color = 2'b00;
		14'h3dbb: color = 2'b00;
		14'h3dbc: color = 2'b10;
		14'h3dbd: color = 2'b11;
		14'h3dbe: color = 2'b11;
		14'h3dbf: color = 2'b11;
		14'h3dc0: color = 2'b10;
		14'h3dc1: color = 2'b11;
		14'h3dc2: color = 2'b11;
		14'h3dc3: color = 2'b10;
		14'h3dc4: color = 2'b01;
		14'h3dc5: color = 2'b10;
		14'h3dc6: color = 2'b10;
		14'h3dc7: color = 2'b11;
		14'h3dc8: color = 2'b11;
		14'h3dc9: color = 2'b10;
		14'h3dca: color = 2'b01;
		14'h3dcb: color = 2'b11;
		14'h3dcc: color = 2'b01;
		14'h3dcd: color = 2'b10;
		14'h3dce: color = 2'b11;
		14'h3dcf: color = 2'b11;
		14'h3dd0: color = 2'b11;
		14'h3dd1: color = 2'b11;
		14'h3dd2: color = 2'b11;
		14'h3dd3: color = 2'b01;
		14'h3dd4: color = 2'b01;
		14'h3dd5: color = 2'b00;
		14'h3dd6: color = 2'b00;
		14'h3dd7: color = 2'b00;
		14'h3dd8: color = 2'b00;
		14'h3dd9: color = 2'b00;
		14'h3dda: color = 2'b00;
		14'h3ddb: color = 2'b00;
		14'h3ddc: color = 2'b00;
		14'h3ddd: color = 2'b00;
		14'h3dde: color = 2'b00;
		14'h3ddf: color = 2'b00;
		14'h3de0: color = 2'b00;
		14'h3de1: color = 2'b00;
		14'h3de2: color = 2'b00;
		14'h3de3: color = 2'b00;
		14'h3de4: color = 2'b00;
		14'h3de5: color = 2'b00;
		14'h3de6: color = 2'b00;
		14'h3de7: color = 2'b00;
		14'h3de8: color = 2'b00;
		14'h3de9: color = 2'b00;
		14'h3dea: color = 2'b00;
		14'h3deb: color = 2'b00;
		14'h3dec: color = 2'b00;
		14'h3ded: color = 2'b00;
		14'h3dee: color = 2'b00;
		14'h3def: color = 2'b00;
		14'h3df0: color = 2'b00;
		14'h3df1: color = 2'b00;
		14'h3df2: color = 2'b00;
		14'h3df3: color = 2'b00;
		14'h3df4: color = 2'b00;
		14'h3df5: color = 2'b00;
		14'h3df6: color = 2'b00;
		14'h3df7: color = 2'b00;
		14'h3df8: color = 2'b00;
		14'h3df9: color = 2'b00;
		14'h3dfa: color = 2'b01;
		14'h3dfb: color = 2'b11;
		14'h3dfc: color = 2'b11;
		14'h3dfd: color = 2'b11;
		14'h3dfe: color = 2'b11;
		14'h3dff: color = 2'b11;
		14'h3e00: color = 2'b01;
		14'h3e01: color = 2'b00;
		14'h3e02: color = 2'b00;
		14'h3e03: color = 2'b00;
		14'h3e04: color = 2'b00;
		14'h3e05: color = 2'b00;
		14'h3e06: color = 2'b00;
		14'h3e07: color = 2'b00;
		14'h3e08: color = 2'b00;
		14'h3e09: color = 2'b00;
		14'h3e0a: color = 2'b00;
		14'h3e0b: color = 2'b00;
		14'h3e0c: color = 2'b00;
		14'h3e0d: color = 2'b00;
		14'h3e0e: color = 2'b00;
		14'h3e0f: color = 2'b00;
		14'h3e10: color = 2'b00;
		14'h3e11: color = 2'b00;
		14'h3e12: color = 2'b00;
		14'h3e13: color = 2'b00;
		14'h3e14: color = 2'b00;
		14'h3e15: color = 2'b00;
		14'h3e16: color = 2'b00;
		14'h3e17: color = 2'b00;
		14'h3e18: color = 2'b00;
		14'h3e19: color = 2'b00;
		14'h3e1a: color = 2'b00;
		14'h3e1b: color = 2'b00;
		14'h3e1c: color = 2'b00;
		14'h3e1d: color = 2'b00;
		14'h3e1e: color = 2'b00;
		14'h3e1f: color = 2'b00;
		14'h3e20: color = 2'b00;
		14'h3e21: color = 2'b00;
		14'h3e22: color = 2'b00;
		14'h3e23: color = 2'b00;
		14'h3e24: color = 2'b00;
		14'h3e25: color = 2'b00;
		14'h3e26: color = 2'b00;
		14'h3e27: color = 2'b00;
		14'h3e28: color = 2'b00;
		14'h3e29: color = 2'b00;
		14'h3e2a: color = 2'b00;
		14'h3e2b: color = 2'b00;
		14'h3e2c: color = 2'b00;
		14'h3e2d: color = 2'b00;
		14'h3e2e: color = 2'b00;
		14'h3e2f: color = 2'b00;
		14'h3e30: color = 2'b00;
		14'h3e31: color = 2'b00;
		14'h3e32: color = 2'b00;
		14'h3e33: color = 2'b00;
		14'h3e34: color = 2'b00;
		14'h3e35: color = 2'b00;
		14'h3e36: color = 2'b00;
		14'h3e37: color = 2'b00;
		14'h3e38: color = 2'b00;
		14'h3e39: color = 2'b00;
		14'h3e3a: color = 2'b00;
		14'h3e3b: color = 2'b00;
		14'h3e3c: color = 2'b00;
		14'h3e3d: color = 2'b11;
		14'h3e3e: color = 2'b11;
		14'h3e3f: color = 2'b11;
		14'h3e40: color = 2'b10;
		14'h3e41: color = 2'b11;
		14'h3e42: color = 2'b10;
		14'h3e43: color = 2'b10;
		14'h3e44: color = 2'b01;
		14'h3e45: color = 2'b10;
		14'h3e46: color = 2'b11;
		14'h3e47: color = 2'b10;
		14'h3e48: color = 2'b10;
		14'h3e49: color = 2'b01;
		14'h3e4a: color = 2'b01;
		14'h3e4b: color = 2'b11;
		14'h3e4c: color = 2'b01;
		14'h3e4d: color = 2'b10;
		14'h3e4e: color = 2'b10;
		14'h3e4f: color = 2'b11;
		14'h3e50: color = 2'b11;
		14'h3e51: color = 2'b11;
		14'h3e52: color = 2'b11;
		14'h3e53: color = 2'b10;
		14'h3e54: color = 2'b00;
		14'h3e55: color = 2'b00;
		14'h3e56: color = 2'b00;
		14'h3e57: color = 2'b00;
		14'h3e58: color = 2'b00;
		14'h3e59: color = 2'b00;
		14'h3e5a: color = 2'b00;
		14'h3e5b: color = 2'b00;
		14'h3e5c: color = 2'b00;
		14'h3e5d: color = 2'b00;
		14'h3e5e: color = 2'b00;
		14'h3e5f: color = 2'b00;
		14'h3e60: color = 2'b00;
		14'h3e61: color = 2'b00;
		14'h3e62: color = 2'b00;
		14'h3e63: color = 2'b00;
		14'h3e64: color = 2'b00;
		14'h3e65: color = 2'b00;
		14'h3e66: color = 2'b00;
		14'h3e67: color = 2'b00;
		14'h3e68: color = 2'b00;
		14'h3e69: color = 2'b00;
		14'h3e6a: color = 2'b00;
		14'h3e6b: color = 2'b00;
		14'h3e6c: color = 2'b00;
		14'h3e6d: color = 2'b00;
		14'h3e6e: color = 2'b00;
		14'h3e6f: color = 2'b00;
		14'h3e70: color = 2'b00;
		14'h3e71: color = 2'b00;
		14'h3e72: color = 2'b00;
		14'h3e73: color = 2'b00;
		14'h3e74: color = 2'b00;
		14'h3e75: color = 2'b00;
		14'h3e76: color = 2'b00;
		14'h3e77: color = 2'b00;
		14'h3e78: color = 2'b00;
		14'h3e79: color = 2'b00;
		14'h3e7a: color = 2'b00;
		14'h3e7b: color = 2'b11;
		14'h3e7c: color = 2'b11;
		14'h3e7d: color = 2'b11;
		14'h3e7e: color = 2'b11;
		14'h3e7f: color = 2'b11;
		14'h3e80: color = 2'b01;
		14'h3e81: color = 2'b00;
		14'h3e82: color = 2'b01;
		14'h3e83: color = 2'b00;
		14'h3e84: color = 2'b00;
		14'h3e85: color = 2'b00;
		14'h3e86: color = 2'b00;
		14'h3e87: color = 2'b00;
		14'h3e88: color = 2'b00;
		14'h3e89: color = 2'b00;
		14'h3e8a: color = 2'b00;
		14'h3e8b: color = 2'b00;
		14'h3e8c: color = 2'b00;
		14'h3e8d: color = 2'b00;
		14'h3e8e: color = 2'b00;
		14'h3e8f: color = 2'b00;
		14'h3e90: color = 2'b00;
		14'h3e91: color = 2'b00;
		14'h3e92: color = 2'b00;
		14'h3e93: color = 2'b00;
		14'h3e94: color = 2'b00;
		14'h3e95: color = 2'b00;
		14'h3e96: color = 2'b00;
		14'h3e97: color = 2'b00;
		14'h3e98: color = 2'b00;
		14'h3e99: color = 2'b00;
		14'h3e9a: color = 2'b00;
		14'h3e9b: color = 2'b00;
		14'h3e9c: color = 2'b00;
		14'h3e9d: color = 2'b00;
		14'h3e9e: color = 2'b00;
		14'h3e9f: color = 2'b00;
		14'h3ea0: color = 2'b00;
		14'h3ea1: color = 2'b00;
		14'h3ea2: color = 2'b00;
		14'h3ea3: color = 2'b00;
		14'h3ea4: color = 2'b00;
		14'h3ea5: color = 2'b00;
		14'h3ea6: color = 2'b00;
		14'h3ea7: color = 2'b00;
		14'h3ea8: color = 2'b00;
		14'h3ea9: color = 2'b00;
		14'h3eaa: color = 2'b00;
		14'h3eab: color = 2'b00;
		14'h3eac: color = 2'b00;
		14'h3ead: color = 2'b00;
		14'h3eae: color = 2'b00;
		14'h3eaf: color = 2'b00;
		14'h3eb0: color = 2'b00;
		14'h3eb1: color = 2'b00;
		14'h3eb2: color = 2'b00;
		14'h3eb3: color = 2'b00;
		14'h3eb4: color = 2'b00;
		14'h3eb5: color = 2'b00;
		14'h3eb6: color = 2'b00;
		14'h3eb7: color = 2'b00;
		14'h3eb8: color = 2'b00;
		14'h3eb9: color = 2'b00;
		14'h3eba: color = 2'b00;
		14'h3ebb: color = 2'b00;
		14'h3ebc: color = 2'b00;
		14'h3ebd: color = 2'b10;
		14'h3ebe: color = 2'b11;
		14'h3ebf: color = 2'b10;
		14'h3ec0: color = 2'b10;
		14'h3ec1: color = 2'b11;
		14'h3ec2: color = 2'b10;
		14'h3ec3: color = 2'b01;
		14'h3ec4: color = 2'b10;
		14'h3ec5: color = 2'b10;
		14'h3ec6: color = 2'b10;
		14'h3ec7: color = 2'b10;
		14'h3ec8: color = 2'b10;
		14'h3ec9: color = 2'b01;
		14'h3eca: color = 2'b01;
		14'h3ecb: color = 2'b11;
		14'h3ecc: color = 2'b01;
		14'h3ecd: color = 2'b01;
		14'h3ece: color = 2'b11;
		14'h3ecf: color = 2'b11;
		14'h3ed0: color = 2'b11;
		14'h3ed1: color = 2'b10;
		14'h3ed2: color = 2'b11;
		14'h3ed3: color = 2'b10;
		14'h3ed4: color = 2'b01;
		14'h3ed5: color = 2'b00;
		14'h3ed6: color = 2'b00;
		14'h3ed7: color = 2'b00;
		14'h3ed8: color = 2'b00;
		14'h3ed9: color = 2'b00;
		14'h3eda: color = 2'b00;
		14'h3edb: color = 2'b00;
		14'h3edc: color = 2'b00;
		14'h3edd: color = 2'b00;
		14'h3ede: color = 2'b00;
		14'h3edf: color = 2'b00;
		14'h3ee0: color = 2'b00;
		14'h3ee1: color = 2'b00;
		14'h3ee2: color = 2'b00;
		14'h3ee3: color = 2'b00;
		14'h3ee4: color = 2'b00;
		14'h3ee5: color = 2'b00;
		14'h3ee6: color = 2'b00;
		14'h3ee7: color = 2'b00;
		14'h3ee8: color = 2'b00;
		14'h3ee9: color = 2'b00;
		14'h3eea: color = 2'b00;
		14'h3eeb: color = 2'b00;
		14'h3eec: color = 2'b00;
		14'h3eed: color = 2'b00;
		14'h3eee: color = 2'b00;
		14'h3eef: color = 2'b00;
		14'h3ef0: color = 2'b00;
		14'h3ef1: color = 2'b00;
		14'h3ef2: color = 2'b00;
		14'h3ef3: color = 2'b00;
		14'h3ef4: color = 2'b00;
		14'h3ef5: color = 2'b00;
		14'h3ef6: color = 2'b00;
		14'h3ef7: color = 2'b00;
		14'h3ef8: color = 2'b00;
		14'h3ef9: color = 2'b00;
		14'h3efa: color = 2'b00;
		14'h3efb: color = 2'b11;
		14'h3efc: color = 2'b11;
		14'h3efd: color = 2'b11;
		14'h3efe: color = 2'b11;
		14'h3eff: color = 2'b11;
		14'h3f00: color = 2'b01;
		14'h3f01: color = 2'b00;
		14'h3f02: color = 2'b01;
		14'h3f03: color = 2'b00;
		14'h3f04: color = 2'b00;
		14'h3f05: color = 2'b00;
		14'h3f06: color = 2'b00;
		14'h3f07: color = 2'b00;
		14'h3f08: color = 2'b00;
		14'h3f09: color = 2'b00;
		14'h3f0a: color = 2'b00;
		14'h3f0b: color = 2'b00;
		14'h3f0c: color = 2'b00;
		14'h3f0d: color = 2'b00;
		14'h3f0e: color = 2'b00;
		14'h3f0f: color = 2'b00;
		14'h3f10: color = 2'b00;
		14'h3f11: color = 2'b00;
		14'h3f12: color = 2'b00;
		14'h3f13: color = 2'b00;
		14'h3f14: color = 2'b00;
		14'h3f15: color = 2'b00;
		14'h3f16: color = 2'b00;
		14'h3f17: color = 2'b00;
		14'h3f18: color = 2'b00;
		14'h3f19: color = 2'b00;
		14'h3f1a: color = 2'b00;
		14'h3f1b: color = 2'b00;
		14'h3f1c: color = 2'b00;
		14'h3f1d: color = 2'b00;
		14'h3f1e: color = 2'b00;
		14'h3f1f: color = 2'b00;
		14'h3f20: color = 2'b00;
		14'h3f21: color = 2'b00;
		14'h3f22: color = 2'b00;
		14'h3f23: color = 2'b00;
		14'h3f24: color = 2'b00;
		14'h3f25: color = 2'b00;
		14'h3f26: color = 2'b00;
		14'h3f27: color = 2'b00;
		14'h3f28: color = 2'b00;
		14'h3f29: color = 2'b00;
		14'h3f2a: color = 2'b00;
		14'h3f2b: color = 2'b00;
		14'h3f2c: color = 2'b00;
		14'h3f2d: color = 2'b00;
		14'h3f2e: color = 2'b00;
		14'h3f2f: color = 2'b00;
		14'h3f30: color = 2'b00;
		14'h3f31: color = 2'b00;
		14'h3f32: color = 2'b00;
		14'h3f33: color = 2'b00;
		14'h3f34: color = 2'b00;
		14'h3f35: color = 2'b00;
		14'h3f36: color = 2'b00;
		14'h3f37: color = 2'b00;
		14'h3f38: color = 2'b00;
		14'h3f39: color = 2'b00;
		14'h3f3a: color = 2'b00;
		14'h3f3b: color = 2'b00;
		14'h3f3c: color = 2'b00;
		14'h3f3d: color = 2'b01;
		14'h3f3e: color = 2'b11;
		14'h3f3f: color = 2'b11;
		14'h3f40: color = 2'b10;
		14'h3f41: color = 2'b10;
		14'h3f42: color = 2'b01;
		14'h3f43: color = 2'b01;
		14'h3f44: color = 2'b10;
		14'h3f45: color = 2'b10;
		14'h3f46: color = 2'b10;
		14'h3f47: color = 2'b10;
		14'h3f48: color = 2'b10;
		14'h3f49: color = 2'b01;
		14'h3f4a: color = 2'b01;
		14'h3f4b: color = 2'b10;
		14'h3f4c: color = 2'b10;
		14'h3f4d: color = 2'b01;
		14'h3f4e: color = 2'b10;
		14'h3f4f: color = 2'b10;
		14'h3f50: color = 2'b11;
		14'h3f51: color = 2'b11;
		14'h3f52: color = 2'b11;
		14'h3f53: color = 2'b11;
		14'h3f54: color = 2'b10;
		14'h3f55: color = 2'b00;
		14'h3f56: color = 2'b00;
		14'h3f57: color = 2'b00;
		14'h3f58: color = 2'b00;
		14'h3f59: color = 2'b00;
		14'h3f5a: color = 2'b00;
		14'h3f5b: color = 2'b00;
		14'h3f5c: color = 2'b00;
		14'h3f5d: color = 2'b00;
		14'h3f5e: color = 2'b00;
		14'h3f5f: color = 2'b00;
		14'h3f60: color = 2'b00;
		14'h3f61: color = 2'b00;
		14'h3f62: color = 2'b00;
		14'h3f63: color = 2'b00;
		14'h3f64: color = 2'b00;
		14'h3f65: color = 2'b00;
		14'h3f66: color = 2'b00;
		14'h3f67: color = 2'b00;
		14'h3f68: color = 2'b00;
		14'h3f69: color = 2'b00;
		14'h3f6a: color = 2'b00;
		14'h3f6b: color = 2'b00;
		14'h3f6c: color = 2'b00;
		14'h3f6d: color = 2'b00;
		14'h3f6e: color = 2'b00;
		14'h3f6f: color = 2'b00;
		14'h3f70: color = 2'b00;
		14'h3f71: color = 2'b00;
		14'h3f72: color = 2'b00;
		14'h3f73: color = 2'b00;
		14'h3f74: color = 2'b00;
		14'h3f75: color = 2'b00;
		14'h3f76: color = 2'b00;
		14'h3f77: color = 2'b00;
		14'h3f78: color = 2'b00;
		14'h3f79: color = 2'b00;
		14'h3f7a: color = 2'b00;
		14'h3f7b: color = 2'b11;
		14'h3f7c: color = 2'b11;
		14'h3f7d: color = 2'b11;
		14'h3f7e: color = 2'b11;
		14'h3f7f: color = 2'b11;
		14'h3f80: color = 2'b00;
		14'h3f81: color = 2'b00;
		14'h3f82: color = 2'b00;
		14'h3f83: color = 2'b00;
		14'h3f84: color = 2'b00;
		14'h3f85: color = 2'b01;
		14'h3f86: color = 2'b00;
		14'h3f87: color = 2'b00;
		14'h3f88: color = 2'b00;
		14'h3f89: color = 2'b00;
		14'h3f8a: color = 2'b00;
		14'h3f8b: color = 2'b00;
		14'h3f8c: color = 2'b00;
		14'h3f8d: color = 2'b00;
		14'h3f8e: color = 2'b00;
		14'h3f8f: color = 2'b00;
		14'h3f90: color = 2'b00;
		14'h3f91: color = 2'b00;
		14'h3f92: color = 2'b00;
		14'h3f93: color = 2'b00;
		14'h3f94: color = 2'b00;
		14'h3f95: color = 2'b00;
		14'h3f96: color = 2'b00;
		14'h3f97: color = 2'b00;
		14'h3f98: color = 2'b00;
		14'h3f99: color = 2'b00;
		14'h3f9a: color = 2'b00;
		14'h3f9b: color = 2'b00;
		14'h3f9c: color = 2'b00;
		14'h3f9d: color = 2'b00;
		14'h3f9e: color = 2'b00;
		14'h3f9f: color = 2'b00;
		14'h3fa0: color = 2'b00;
		14'h3fa1: color = 2'b00;
		14'h3fa2: color = 2'b00;
		14'h3fa3: color = 2'b00;
		14'h3fa4: color = 2'b00;
		14'h3fa5: color = 2'b00;
		14'h3fa6: color = 2'b00;
		14'h3fa7: color = 2'b00;
		14'h3fa8: color = 2'b00;
		14'h3fa9: color = 2'b00;
		14'h3faa: color = 2'b00;
		14'h3fab: color = 2'b00;
		14'h3fac: color = 2'b00;
		14'h3fad: color = 2'b00;
		14'h3fae: color = 2'b00;
		14'h3faf: color = 2'b00;
		14'h3fb0: color = 2'b00;
		14'h3fb1: color = 2'b00;
		14'h3fb2: color = 2'b00;
		14'h3fb3: color = 2'b00;
		14'h3fb4: color = 2'b00;
		14'h3fb5: color = 2'b00;
		14'h3fb6: color = 2'b00;
		14'h3fb7: color = 2'b00;
		14'h3fb8: color = 2'b00;
		14'h3fb9: color = 2'b00;
		14'h3fba: color = 2'b00;
		14'h3fbb: color = 2'b00;
		14'h3fbc: color = 2'b00;
		14'h3fbd: color = 2'b00;
		14'h3fbe: color = 2'b11;
		14'h3fbf: color = 2'b11;
		14'h3fc0: color = 2'b10;
		14'h3fc1: color = 2'b10;
		14'h3fc2: color = 2'b01;
		14'h3fc3: color = 2'b10;
		14'h3fc4: color = 2'b10;
		14'h3fc5: color = 2'b10;
		14'h3fc6: color = 2'b10;
		14'h3fc7: color = 2'b01;
		14'h3fc8: color = 2'b01;
		14'h3fc9: color = 2'b10;
		14'h3fca: color = 2'b10;
		14'h3fcb: color = 2'b11;
		14'h3fcc: color = 2'b10;
		14'h3fcd: color = 2'b10;
		14'h3fce: color = 2'b10;
		14'h3fcf: color = 2'b10;
		14'h3fd0: color = 2'b11;
		14'h3fd1: color = 2'b11;
		14'h3fd2: color = 2'b11;
		14'h3fd3: color = 2'b11;
		14'h3fd4: color = 2'b10;
		14'h3fd5: color = 2'b01;
		14'h3fd6: color = 2'b00;
		14'h3fd7: color = 2'b00;
		14'h3fd8: color = 2'b00;
		14'h3fd9: color = 2'b00;
		14'h3fda: color = 2'b00;
		14'h3fdb: color = 2'b00;
		14'h3fdc: color = 2'b00;
		14'h3fdd: color = 2'b00;
		14'h3fde: color = 2'b00;
		14'h3fdf: color = 2'b00;
		14'h3fe0: color = 2'b00;
		14'h3fe1: color = 2'b00;
		14'h3fe2: color = 2'b00;
		14'h3fe3: color = 2'b00;
		14'h3fe4: color = 2'b00;
		14'h3fe5: color = 2'b00;
		14'h3fe6: color = 2'b00;
		14'h3fe7: color = 2'b00;
		14'h3fe8: color = 2'b00;
		14'h3fe9: color = 2'b00;
		14'h3fea: color = 2'b00;
		14'h3feb: color = 2'b00;
		14'h3fec: color = 2'b00;
		14'h3fed: color = 2'b00;
		14'h3fee: color = 2'b00;
		14'h3fef: color = 2'b00;
		14'h3ff0: color = 2'b00;
		14'h3ff1: color = 2'b00;
		14'h3ff2: color = 2'b00;
		14'h3ff3: color = 2'b00;
		14'h3ff4: color = 2'b00;
		14'h3ff5: color = 2'b00;
		14'h3ff6: color = 2'b00;
		14'h3ff7: color = 2'b00;
		14'h3ff8: color = 2'b00;
		14'h3ff9: color = 2'b00;
		14'h3ffa: color = 2'b00;
		14'h3ffb: color = 2'b11;
		14'h3ffc: color = 2'b11;
		14'h3ffd: color = 2'b11;
		14'h3ffe: color = 2'b11;
		14'h3fff: color = 2'b11;
	endcase
end
endmodule
