module Computer
(
   input            clock, 
   input      [7:0] x,
   input      [7:0] y, 
   input      [7:0] loc_x, 
   input      [7:0] loc_y, 
   output reg       on,
   output reg [1:0] color
);

   localparam WIDTH = 8'd32,
              HEIGHT = 8'd64;

   // Buffer the scan coordinates to synchronize
   // with the ROM data output
   always @( posedge clock ) begin
    on <= (x >= loc_x && x <= (loc_x+(WIDTH-1)))
          && (y >= loc_y && y <= (loc_y+(HEIGHT-1)));
   end

   reg [10:0] addr;
   always @( posedge clock )
      addr <= {y[5:0]-loc_y[5:0],x[4:0]-loc_x[4:0]};

always @(*) begin
   case( addr )
      11'h000: color = 2'b11;
      11'h001: color = 2'b11;
      11'h002: color = 2'b11;
      11'h003: color = 2'b11;
      11'h004: color = 2'b11;
      11'h005: color = 2'b11;
      11'h006: color = 2'b00;
      11'h007: color = 2'b00;
      11'h008: color = 2'b00;
      11'h009: color = 2'b00;
      11'h00a: color = 2'b00;
      11'h00b: color = 2'b00;
      11'h00c: color = 2'b00;
      11'h00d: color = 2'b00;
      11'h00e: color = 2'b00;
      11'h00f: color = 2'b00;
      11'h010: color = 2'b00;
      11'h011: color = 2'b00;
      11'h012: color = 2'b00;
      11'h013: color = 2'b00;
      11'h014: color = 2'b00;
      11'h015: color = 2'b00;
      11'h016: color = 2'b00;
      11'h017: color = 2'b00;
      11'h018: color = 2'b00;
      11'h019: color = 2'b00;
      11'h01a: color = 2'b11;
      11'h01b: color = 2'b11;
      11'h01c: color = 2'b11;
      11'h01d: color = 2'b11;
      11'h01e: color = 2'b11;
      11'h01f: color = 2'b11;
      11'h020: color = 2'b11;
      11'h021: color = 2'b11;
      11'h022: color = 2'b11;
      11'h023: color = 2'b11;
      11'h024: color = 2'b11;
      11'h025: color = 2'b11;
      11'h026: color = 2'b00;
      11'h027: color = 2'b00;
      11'h028: color = 2'b00;
      11'h029: color = 2'b00;
      11'h02a: color = 2'b00;
      11'h02b: color = 2'b00;
      11'h02c: color = 2'b00;
      11'h02d: color = 2'b00;
      11'h02e: color = 2'b00;
      11'h02f: color = 2'b00;
      11'h030: color = 2'b00;
      11'h031: color = 2'b00;
      11'h032: color = 2'b00;
      11'h033: color = 2'b00;
      11'h034: color = 2'b00;
      11'h035: color = 2'b00;
      11'h036: color = 2'b00;
      11'h037: color = 2'b00;
      11'h038: color = 2'b00;
      11'h039: color = 2'b00;
      11'h03a: color = 2'b11;
      11'h03b: color = 2'b11;
      11'h03c: color = 2'b11;
      11'h03d: color = 2'b11;
      11'h03e: color = 2'b11;
      11'h03f: color = 2'b11;
      11'h040: color = 2'b11;
      11'h041: color = 2'b11;
      11'h042: color = 2'b11;
      11'h043: color = 2'b11;
      11'h044: color = 2'b00;
      11'h045: color = 2'b00;
      11'h046: color = 2'b11;
      11'h047: color = 2'b11;
      11'h048: color = 2'b11;
      11'h049: color = 2'b11;
      11'h04a: color = 2'b11;
      11'h04b: color = 2'b11;
      11'h04c: color = 2'b11;
      11'h04d: color = 2'b11;
      11'h04e: color = 2'b11;
      11'h04f: color = 2'b11;
      11'h050: color = 2'b11;
      11'h051: color = 2'b11;
      11'h052: color = 2'b11;
      11'h053: color = 2'b11;
      11'h054: color = 2'b11;
      11'h055: color = 2'b11;
      11'h056: color = 2'b11;
      11'h057: color = 2'b11;
      11'h058: color = 2'b11;
      11'h059: color = 2'b11;
      11'h05a: color = 2'b00;
      11'h05b: color = 2'b00;
      11'h05c: color = 2'b11;
      11'h05d: color = 2'b11;
      11'h05e: color = 2'b11;
      11'h05f: color = 2'b11;
      11'h060: color = 2'b11;
      11'h061: color = 2'b11;
      11'h062: color = 2'b11;
      11'h063: color = 2'b11;
      11'h064: color = 2'b00;
      11'h065: color = 2'b00;
      11'h066: color = 2'b11;
      11'h067: color = 2'b11;
      11'h068: color = 2'b11;
      11'h069: color = 2'b11;
      11'h06a: color = 2'b11;
      11'h06b: color = 2'b11;
      11'h06c: color = 2'b11;
      11'h06d: color = 2'b11;
      11'h06e: color = 2'b11;
      11'h06f: color = 2'b11;
      11'h070: color = 2'b11;
      11'h071: color = 2'b11;
      11'h072: color = 2'b11;
      11'h073: color = 2'b11;
      11'h074: color = 2'b11;
      11'h075: color = 2'b11;
      11'h076: color = 2'b11;
      11'h077: color = 2'b11;
      11'h078: color = 2'b11;
      11'h079: color = 2'b11;
      11'h07a: color = 2'b00;
      11'h07b: color = 2'b00;
      11'h07c: color = 2'b11;
      11'h07d: color = 2'b11;
      11'h07e: color = 2'b11;
      11'h07f: color = 2'b11;
      11'h080: color = 2'b11;
      11'h081: color = 2'b11;
      11'h082: color = 2'b11;
      11'h083: color = 2'b11;
      11'h084: color = 2'b00;
      11'h085: color = 2'b00;
      11'h086: color = 2'b11;
      11'h087: color = 2'b11;
      11'h088: color = 2'b11;
      11'h089: color = 2'b11;
      11'h08a: color = 2'b11;
      11'h08b: color = 2'b11;
      11'h08c: color = 2'b11;
      11'h08d: color = 2'b11;
      11'h08e: color = 2'b11;
      11'h08f: color = 2'b11;
      11'h090: color = 2'b11;
      11'h091: color = 2'b11;
      11'h092: color = 2'b11;
      11'h093: color = 2'b11;
      11'h094: color = 2'b11;
      11'h095: color = 2'b11;
      11'h096: color = 2'b11;
      11'h097: color = 2'b11;
      11'h098: color = 2'b11;
      11'h099: color = 2'b11;
      11'h09a: color = 2'b00;
      11'h09b: color = 2'b00;
      11'h09c: color = 2'b11;
      11'h09d: color = 2'b11;
      11'h09e: color = 2'b11;
      11'h09f: color = 2'b11;
      11'h0a0: color = 2'b11;
      11'h0a1: color = 2'b11;
      11'h0a2: color = 2'b11;
      11'h0a3: color = 2'b11;
      11'h0a4: color = 2'b00;
      11'h0a5: color = 2'b00;
      11'h0a6: color = 2'b11;
      11'h0a7: color = 2'b11;
      11'h0a8: color = 2'b11;
      11'h0a9: color = 2'b11;
      11'h0aa: color = 2'b11;
      11'h0ab: color = 2'b11;
      11'h0ac: color = 2'b11;
      11'h0ad: color = 2'b11;
      11'h0ae: color = 2'b11;
      11'h0af: color = 2'b11;
      11'h0b0: color = 2'b11;
      11'h0b1: color = 2'b11;
      11'h0b2: color = 2'b11;
      11'h0b3: color = 2'b11;
      11'h0b4: color = 2'b11;
      11'h0b5: color = 2'b11;
      11'h0b6: color = 2'b11;
      11'h0b7: color = 2'b11;
      11'h0b8: color = 2'b11;
      11'h0b9: color = 2'b11;
      11'h0ba: color = 2'b00;
      11'h0bb: color = 2'b00;
      11'h0bc: color = 2'b11;
      11'h0bd: color = 2'b11;
      11'h0be: color = 2'b11;
      11'h0bf: color = 2'b11;
      11'h0c0: color = 2'b11;
      11'h0c1: color = 2'b11;
      11'h0c2: color = 2'b11;
      11'h0c3: color = 2'b11;
      11'h0c4: color = 2'b00;
      11'h0c5: color = 2'b00;
      11'h0c6: color = 2'b11;
      11'h0c7: color = 2'b11;
      11'h0c8: color = 2'b11;
      11'h0c9: color = 2'b11;
      11'h0ca: color = 2'b11;
      11'h0cb: color = 2'b11;
      11'h0cc: color = 2'b11;
      11'h0cd: color = 2'b11;
      11'h0ce: color = 2'b11;
      11'h0cf: color = 2'b11;
      11'h0d0: color = 2'b11;
      11'h0d1: color = 2'b11;
      11'h0d2: color = 2'b11;
      11'h0d3: color = 2'b11;
      11'h0d4: color = 2'b11;
      11'h0d5: color = 2'b11;
      11'h0d6: color = 2'b11;
      11'h0d7: color = 2'b11;
      11'h0d8: color = 2'b11;
      11'h0d9: color = 2'b11;
      11'h0da: color = 2'b00;
      11'h0db: color = 2'b00;
      11'h0dc: color = 2'b11;
      11'h0dd: color = 2'b11;
      11'h0de: color = 2'b11;
      11'h0df: color = 2'b11;
      11'h0e0: color = 2'b11;
      11'h0e1: color = 2'b11;
      11'h0e2: color = 2'b11;
      11'h0e3: color = 2'b11;
      11'h0e4: color = 2'b00;
      11'h0e5: color = 2'b00;
      11'h0e6: color = 2'b11;
      11'h0e7: color = 2'b11;
      11'h0e8: color = 2'b11;
      11'h0e9: color = 2'b11;
      11'h0ea: color = 2'b11;
      11'h0eb: color = 2'b11;
      11'h0ec: color = 2'b11;
      11'h0ed: color = 2'b11;
      11'h0ee: color = 2'b11;
      11'h0ef: color = 2'b11;
      11'h0f0: color = 2'b11;
      11'h0f1: color = 2'b11;
      11'h0f2: color = 2'b11;
      11'h0f3: color = 2'b11;
      11'h0f4: color = 2'b11;
      11'h0f5: color = 2'b11;
      11'h0f6: color = 2'b11;
      11'h0f7: color = 2'b11;
      11'h0f8: color = 2'b11;
      11'h0f9: color = 2'b11;
      11'h0fa: color = 2'b00;
      11'h0fb: color = 2'b00;
      11'h0fc: color = 2'b11;
      11'h0fd: color = 2'b11;
      11'h0fe: color = 2'b11;
      11'h0ff: color = 2'b11;
      11'h100: color = 2'b11;
      11'h101: color = 2'b11;
      11'h102: color = 2'b11;
      11'h103: color = 2'b11;
      11'h104: color = 2'b00;
      11'h105: color = 2'b00;
      11'h106: color = 2'b10;
      11'h107: color = 2'b10;
      11'h108: color = 2'b10;
      11'h109: color = 2'b10;
      11'h10a: color = 2'b10;
      11'h10b: color = 2'b10;
      11'h10c: color = 2'b10;
      11'h10d: color = 2'b10;
      11'h10e: color = 2'b10;
      11'h10f: color = 2'b10;
      11'h110: color = 2'b10;
      11'h111: color = 2'b10;
      11'h112: color = 2'b10;
      11'h113: color = 2'b10;
      11'h114: color = 2'b10;
      11'h115: color = 2'b10;
      11'h116: color = 2'b10;
      11'h117: color = 2'b10;
      11'h118: color = 2'b10;
      11'h119: color = 2'b10;
      11'h11a: color = 2'b00;
      11'h11b: color = 2'b00;
      11'h11c: color = 2'b11;
      11'h11d: color = 2'b11;
      11'h11e: color = 2'b11;
      11'h11f: color = 2'b11;
      11'h120: color = 2'b11;
      11'h121: color = 2'b11;
      11'h122: color = 2'b11;
      11'h123: color = 2'b11;
      11'h124: color = 2'b00;
      11'h125: color = 2'b00;
      11'h126: color = 2'b10;
      11'h127: color = 2'b10;
      11'h128: color = 2'b10;
      11'h129: color = 2'b10;
      11'h12a: color = 2'b10;
      11'h12b: color = 2'b10;
      11'h12c: color = 2'b10;
      11'h12d: color = 2'b10;
      11'h12e: color = 2'b10;
      11'h12f: color = 2'b10;
      11'h130: color = 2'b10;
      11'h131: color = 2'b10;
      11'h132: color = 2'b10;
      11'h133: color = 2'b10;
      11'h134: color = 2'b10;
      11'h135: color = 2'b10;
      11'h136: color = 2'b10;
      11'h137: color = 2'b10;
      11'h138: color = 2'b10;
      11'h139: color = 2'b10;
      11'h13a: color = 2'b00;
      11'h13b: color = 2'b00;
      11'h13c: color = 2'b11;
      11'h13d: color = 2'b11;
      11'h13e: color = 2'b11;
      11'h13f: color = 2'b11;
      11'h140: color = 2'b11;
      11'h141: color = 2'b11;
      11'h142: color = 2'b11;
      11'h143: color = 2'b11;
      11'h144: color = 2'b00;
      11'h145: color = 2'b00;
      11'h146: color = 2'b10;
      11'h147: color = 2'b10;
      11'h148: color = 2'b00;
      11'h149: color = 2'b00;
      11'h14a: color = 2'b00;
      11'h14b: color = 2'b00;
      11'h14c: color = 2'b00;
      11'h14d: color = 2'b00;
      11'h14e: color = 2'b00;
      11'h14f: color = 2'b00;
      11'h150: color = 2'b00;
      11'h151: color = 2'b00;
      11'h152: color = 2'b00;
      11'h153: color = 2'b00;
      11'h154: color = 2'b00;
      11'h155: color = 2'b00;
      11'h156: color = 2'b00;
      11'h157: color = 2'b00;
      11'h158: color = 2'b10;
      11'h159: color = 2'b10;
      11'h15a: color = 2'b00;
      11'h15b: color = 2'b00;
      11'h15c: color = 2'b11;
      11'h15d: color = 2'b11;
      11'h15e: color = 2'b11;
      11'h15f: color = 2'b11;
      11'h160: color = 2'b11;
      11'h161: color = 2'b11;
      11'h162: color = 2'b11;
      11'h163: color = 2'b11;
      11'h164: color = 2'b00;
      11'h165: color = 2'b00;
      11'h166: color = 2'b10;
      11'h167: color = 2'b10;
      11'h168: color = 2'b00;
      11'h169: color = 2'b00;
      11'h16a: color = 2'b00;
      11'h16b: color = 2'b00;
      11'h16c: color = 2'b00;
      11'h16d: color = 2'b00;
      11'h16e: color = 2'b00;
      11'h16f: color = 2'b00;
      11'h170: color = 2'b00;
      11'h171: color = 2'b00;
      11'h172: color = 2'b00;
      11'h173: color = 2'b00;
      11'h174: color = 2'b00;
      11'h175: color = 2'b00;
      11'h176: color = 2'b00;
      11'h177: color = 2'b00;
      11'h178: color = 2'b10;
      11'h179: color = 2'b10;
      11'h17a: color = 2'b00;
      11'h17b: color = 2'b00;
      11'h17c: color = 2'b11;
      11'h17d: color = 2'b11;
      11'h17e: color = 2'b11;
      11'h17f: color = 2'b11;
      11'h180: color = 2'b00;
      11'h181: color = 2'b00;
      11'h182: color = 2'b00;
      11'h183: color = 2'b00;
      11'h184: color = 2'b00;
      11'h185: color = 2'b00;
      11'h186: color = 2'b10;
      11'h187: color = 2'b10;
      11'h188: color = 2'b00;
      11'h189: color = 2'b00;
      11'h18a: color = 2'b11;
      11'h18b: color = 2'b11;
      11'h18c: color = 2'b01;
      11'h18d: color = 2'b01;
      11'h18e: color = 2'b00;
      11'h18f: color = 2'b00;
      11'h190: color = 2'b00;
      11'h191: color = 2'b00;
      11'h192: color = 2'b00;
      11'h193: color = 2'b00;
      11'h194: color = 2'b00;
      11'h195: color = 2'b00;
      11'h196: color = 2'b00;
      11'h197: color = 2'b00;
      11'h198: color = 2'b10;
      11'h199: color = 2'b10;
      11'h19a: color = 2'b00;
      11'h19b: color = 2'b00;
      11'h19c: color = 2'b00;
      11'h19d: color = 2'b00;
      11'h19e: color = 2'b00;
      11'h19f: color = 2'b00;
      11'h1a0: color = 2'b00;
      11'h1a1: color = 2'b00;
      11'h1a2: color = 2'b00;
      11'h1a3: color = 2'b00;
      11'h1a4: color = 2'b00;
      11'h1a5: color = 2'b00;
      11'h1a6: color = 2'b10;
      11'h1a7: color = 2'b10;
      11'h1a8: color = 2'b00;
      11'h1a9: color = 2'b00;
      11'h1aa: color = 2'b11;
      11'h1ab: color = 2'b11;
      11'h1ac: color = 2'b01;
      11'h1ad: color = 2'b01;
      11'h1ae: color = 2'b00;
      11'h1af: color = 2'b00;
      11'h1b0: color = 2'b00;
      11'h1b1: color = 2'b00;
      11'h1b2: color = 2'b00;
      11'h1b3: color = 2'b00;
      11'h1b4: color = 2'b00;
      11'h1b5: color = 2'b00;
      11'h1b6: color = 2'b00;
      11'h1b7: color = 2'b00;
      11'h1b8: color = 2'b10;
      11'h1b9: color = 2'b10;
      11'h1ba: color = 2'b00;
      11'h1bb: color = 2'b00;
      11'h1bc: color = 2'b00;
      11'h1bd: color = 2'b00;
      11'h1be: color = 2'b00;
      11'h1bf: color = 2'b00;
      11'h1c0: color = 2'b00;
      11'h1c1: color = 2'b00;
      11'h1c2: color = 2'b11;
      11'h1c3: color = 2'b11;
      11'h1c4: color = 2'b00;
      11'h1c5: color = 2'b00;
      11'h1c6: color = 2'b10;
      11'h1c7: color = 2'b10;
      11'h1c8: color = 2'b00;
      11'h1c9: color = 2'b00;
      11'h1ca: color = 2'b00;
      11'h1cb: color = 2'b00;
      11'h1cc: color = 2'b00;
      11'h1cd: color = 2'b00;
      11'h1ce: color = 2'b00;
      11'h1cf: color = 2'b00;
      11'h1d0: color = 2'b00;
      11'h1d1: color = 2'b00;
      11'h1d2: color = 2'b00;
      11'h1d3: color = 2'b00;
      11'h1d4: color = 2'b00;
      11'h1d5: color = 2'b00;
      11'h1d6: color = 2'b00;
      11'h1d7: color = 2'b00;
      11'h1d8: color = 2'b10;
      11'h1d9: color = 2'b10;
      11'h1da: color = 2'b00;
      11'h1db: color = 2'b00;
      11'h1dc: color = 2'b10;
      11'h1dd: color = 2'b10;
      11'h1de: color = 2'b00;
      11'h1df: color = 2'b00;
      11'h1e0: color = 2'b00;
      11'h1e1: color = 2'b00;
      11'h1e2: color = 2'b11;
      11'h1e3: color = 2'b11;
      11'h1e4: color = 2'b00;
      11'h1e5: color = 2'b00;
      11'h1e6: color = 2'b10;
      11'h1e7: color = 2'b10;
      11'h1e8: color = 2'b00;
      11'h1e9: color = 2'b00;
      11'h1ea: color = 2'b00;
      11'h1eb: color = 2'b00;
      11'h1ec: color = 2'b00;
      11'h1ed: color = 2'b00;
      11'h1ee: color = 2'b00;
      11'h1ef: color = 2'b00;
      11'h1f0: color = 2'b00;
      11'h1f1: color = 2'b00;
      11'h1f2: color = 2'b00;
      11'h1f3: color = 2'b00;
      11'h1f4: color = 2'b00;
      11'h1f5: color = 2'b00;
      11'h1f6: color = 2'b00;
      11'h1f7: color = 2'b00;
      11'h1f8: color = 2'b10;
      11'h1f9: color = 2'b10;
      11'h1fa: color = 2'b00;
      11'h1fb: color = 2'b00;
      11'h1fc: color = 2'b10;
      11'h1fd: color = 2'b10;
      11'h1fe: color = 2'b00;
      11'h1ff: color = 2'b00;
      11'h200: color = 2'b00;
      11'h201: color = 2'b00;
      11'h202: color = 2'b11;
      11'h203: color = 2'b11;
      11'h204: color = 2'b00;
      11'h205: color = 2'b00;
      11'h206: color = 2'b10;
      11'h207: color = 2'b10;
      11'h208: color = 2'b00;
      11'h209: color = 2'b00;
      11'h20a: color = 2'b00;
      11'h20b: color = 2'b00;
      11'h20c: color = 2'b00;
      11'h20d: color = 2'b00;
      11'h20e: color = 2'b00;
      11'h20f: color = 2'b00;
      11'h210: color = 2'b00;
      11'h211: color = 2'b00;
      11'h212: color = 2'b00;
      11'h213: color = 2'b00;
      11'h214: color = 2'b00;
      11'h215: color = 2'b00;
      11'h216: color = 2'b00;
      11'h217: color = 2'b00;
      11'h218: color = 2'b10;
      11'h219: color = 2'b10;
      11'h21a: color = 2'b00;
      11'h21b: color = 2'b00;
      11'h21c: color = 2'b01;
      11'h21d: color = 2'b01;
      11'h21e: color = 2'b00;
      11'h21f: color = 2'b00;
      11'h220: color = 2'b00;
      11'h221: color = 2'b00;
      11'h222: color = 2'b11;
      11'h223: color = 2'b11;
      11'h224: color = 2'b00;
      11'h225: color = 2'b00;
      11'h226: color = 2'b10;
      11'h227: color = 2'b10;
      11'h228: color = 2'b00;
      11'h229: color = 2'b00;
      11'h22a: color = 2'b00;
      11'h22b: color = 2'b00;
      11'h22c: color = 2'b00;
      11'h22d: color = 2'b00;
      11'h22e: color = 2'b00;
      11'h22f: color = 2'b00;
      11'h230: color = 2'b00;
      11'h231: color = 2'b00;
      11'h232: color = 2'b00;
      11'h233: color = 2'b00;
      11'h234: color = 2'b00;
      11'h235: color = 2'b00;
      11'h236: color = 2'b00;
      11'h237: color = 2'b00;
      11'h238: color = 2'b10;
      11'h239: color = 2'b10;
      11'h23a: color = 2'b00;
      11'h23b: color = 2'b00;
      11'h23c: color = 2'b01;
      11'h23d: color = 2'b01;
      11'h23e: color = 2'b00;
      11'h23f: color = 2'b00;
      11'h240: color = 2'b00;
      11'h241: color = 2'b00;
      11'h242: color = 2'b11;
      11'h243: color = 2'b11;
      11'h244: color = 2'b00;
      11'h245: color = 2'b00;
      11'h246: color = 2'b10;
      11'h247: color = 2'b10;
      11'h248: color = 2'b00;
      11'h249: color = 2'b00;
      11'h24a: color = 2'b00;
      11'h24b: color = 2'b00;
      11'h24c: color = 2'b00;
      11'h24d: color = 2'b00;
      11'h24e: color = 2'b00;
      11'h24f: color = 2'b00;
      11'h250: color = 2'b00;
      11'h251: color = 2'b00;
      11'h252: color = 2'b00;
      11'h253: color = 2'b00;
      11'h254: color = 2'b00;
      11'h255: color = 2'b00;
      11'h256: color = 2'b00;
      11'h257: color = 2'b00;
      11'h258: color = 2'b10;
      11'h259: color = 2'b10;
      11'h25a: color = 2'b00;
      11'h25b: color = 2'b00;
      11'h25c: color = 2'b01;
      11'h25d: color = 2'b01;
      11'h25e: color = 2'b00;
      11'h25f: color = 2'b00;
      11'h260: color = 2'b00;
      11'h261: color = 2'b00;
      11'h262: color = 2'b11;
      11'h263: color = 2'b11;
      11'h264: color = 2'b00;
      11'h265: color = 2'b00;
      11'h266: color = 2'b10;
      11'h267: color = 2'b10;
      11'h268: color = 2'b00;
      11'h269: color = 2'b00;
      11'h26a: color = 2'b00;
      11'h26b: color = 2'b00;
      11'h26c: color = 2'b00;
      11'h26d: color = 2'b00;
      11'h26e: color = 2'b00;
      11'h26f: color = 2'b00;
      11'h270: color = 2'b00;
      11'h271: color = 2'b00;
      11'h272: color = 2'b00;
      11'h273: color = 2'b00;
      11'h274: color = 2'b00;
      11'h275: color = 2'b00;
      11'h276: color = 2'b00;
      11'h277: color = 2'b00;
      11'h278: color = 2'b10;
      11'h279: color = 2'b10;
      11'h27a: color = 2'b00;
      11'h27b: color = 2'b00;
      11'h27c: color = 2'b01;
      11'h27d: color = 2'b01;
      11'h27e: color = 2'b00;
      11'h27f: color = 2'b00;
      11'h280: color = 2'b00;
      11'h281: color = 2'b00;
      11'h282: color = 2'b11;
      11'h283: color = 2'b11;
      11'h284: color = 2'b00;
      11'h285: color = 2'b00;
      11'h286: color = 2'b10;
      11'h287: color = 2'b10;
      11'h288: color = 2'b10;
      11'h289: color = 2'b10;
      11'h28a: color = 2'b10;
      11'h28b: color = 2'b10;
      11'h28c: color = 2'b10;
      11'h28d: color = 2'b10;
      11'h28e: color = 2'b10;
      11'h28f: color = 2'b10;
      11'h290: color = 2'b10;
      11'h291: color = 2'b10;
      11'h292: color = 2'b10;
      11'h293: color = 2'b10;
      11'h294: color = 2'b10;
      11'h295: color = 2'b10;
      11'h296: color = 2'b10;
      11'h297: color = 2'b10;
      11'h298: color = 2'b10;
      11'h299: color = 2'b10;
      11'h29a: color = 2'b00;
      11'h29b: color = 2'b00;
      11'h29c: color = 2'b01;
      11'h29d: color = 2'b01;
      11'h29e: color = 2'b00;
      11'h29f: color = 2'b00;
      11'h2a0: color = 2'b00;
      11'h2a1: color = 2'b00;
      11'h2a2: color = 2'b11;
      11'h2a3: color = 2'b11;
      11'h2a4: color = 2'b00;
      11'h2a5: color = 2'b00;
      11'h2a6: color = 2'b10;
      11'h2a7: color = 2'b10;
      11'h2a8: color = 2'b10;
      11'h2a9: color = 2'b10;
      11'h2aa: color = 2'b10;
      11'h2ab: color = 2'b10;
      11'h2ac: color = 2'b10;
      11'h2ad: color = 2'b10;
      11'h2ae: color = 2'b10;
      11'h2af: color = 2'b10;
      11'h2b0: color = 2'b10;
      11'h2b1: color = 2'b10;
      11'h2b2: color = 2'b10;
      11'h2b3: color = 2'b10;
      11'h2b4: color = 2'b10;
      11'h2b5: color = 2'b10;
      11'h2b6: color = 2'b10;
      11'h2b7: color = 2'b10;
      11'h2b8: color = 2'b10;
      11'h2b9: color = 2'b10;
      11'h2ba: color = 2'b00;
      11'h2bb: color = 2'b00;
      11'h2bc: color = 2'b01;
      11'h2bd: color = 2'b01;
      11'h2be: color = 2'b00;
      11'h2bf: color = 2'b00;
      11'h2c0: color = 2'b00;
      11'h2c1: color = 2'b00;
      11'h2c2: color = 2'b11;
      11'h2c3: color = 2'b11;
      11'h2c4: color = 2'b00;
      11'h2c5: color = 2'b00;
      11'h2c6: color = 2'b01;
      11'h2c7: color = 2'b01;
      11'h2c8: color = 2'b01;
      11'h2c9: color = 2'b01;
      11'h2ca: color = 2'b01;
      11'h2cb: color = 2'b01;
      11'h2cc: color = 2'b01;
      11'h2cd: color = 2'b01;
      11'h2ce: color = 2'b01;
      11'h2cf: color = 2'b01;
      11'h2d0: color = 2'b00;
      11'h2d1: color = 2'b00;
      11'h2d2: color = 2'b00;
      11'h2d3: color = 2'b00;
      11'h2d4: color = 2'b00;
      11'h2d5: color = 2'b00;
      11'h2d6: color = 2'b00;
      11'h2d7: color = 2'b00;
      11'h2d8: color = 2'b01;
      11'h2d9: color = 2'b01;
      11'h2da: color = 2'b00;
      11'h2db: color = 2'b00;
      11'h2dc: color = 2'b01;
      11'h2dd: color = 2'b01;
      11'h2de: color = 2'b00;
      11'h2df: color = 2'b00;
      11'h2e0: color = 2'b00;
      11'h2e1: color = 2'b00;
      11'h2e2: color = 2'b11;
      11'h2e3: color = 2'b11;
      11'h2e4: color = 2'b00;
      11'h2e5: color = 2'b00;
      11'h2e6: color = 2'b01;
      11'h2e7: color = 2'b01;
      11'h2e8: color = 2'b01;
      11'h2e9: color = 2'b01;
      11'h2ea: color = 2'b01;
      11'h2eb: color = 2'b01;
      11'h2ec: color = 2'b01;
      11'h2ed: color = 2'b01;
      11'h2ee: color = 2'b01;
      11'h2ef: color = 2'b01;
      11'h2f0: color = 2'b00;
      11'h2f1: color = 2'b00;
      11'h2f2: color = 2'b00;
      11'h2f3: color = 2'b00;
      11'h2f4: color = 2'b00;
      11'h2f5: color = 2'b00;
      11'h2f6: color = 2'b00;
      11'h2f7: color = 2'b00;
      11'h2f8: color = 2'b01;
      11'h2f9: color = 2'b01;
      11'h2fa: color = 2'b00;
      11'h2fb: color = 2'b00;
      11'h2fc: color = 2'b01;
      11'h2fd: color = 2'b01;
      11'h2fe: color = 2'b00;
      11'h2ff: color = 2'b00;
      11'h300: color = 2'b00;
      11'h301: color = 2'b00;
      11'h302: color = 2'b11;
      11'h303: color = 2'b11;
      11'h304: color = 2'b00;
      11'h305: color = 2'b00;
      11'h306: color = 2'b10;
      11'h307: color = 2'b10;
      11'h308: color = 2'b10;
      11'h309: color = 2'b10;
      11'h30a: color = 2'b10;
      11'h30b: color = 2'b10;
      11'h30c: color = 2'b10;
      11'h30d: color = 2'b10;
      11'h30e: color = 2'b10;
      11'h30f: color = 2'b10;
      11'h310: color = 2'b10;
      11'h311: color = 2'b10;
      11'h312: color = 2'b10;
      11'h313: color = 2'b10;
      11'h314: color = 2'b10;
      11'h315: color = 2'b10;
      11'h316: color = 2'b10;
      11'h317: color = 2'b10;
      11'h318: color = 2'b10;
      11'h319: color = 2'b10;
      11'h31a: color = 2'b00;
      11'h31b: color = 2'b00;
      11'h31c: color = 2'b01;
      11'h31d: color = 2'b01;
      11'h31e: color = 2'b00;
      11'h31f: color = 2'b00;
      11'h320: color = 2'b00;
      11'h321: color = 2'b00;
      11'h322: color = 2'b11;
      11'h323: color = 2'b11;
      11'h324: color = 2'b00;
      11'h325: color = 2'b00;
      11'h326: color = 2'b10;
      11'h327: color = 2'b10;
      11'h328: color = 2'b10;
      11'h329: color = 2'b10;
      11'h32a: color = 2'b10;
      11'h32b: color = 2'b10;
      11'h32c: color = 2'b10;
      11'h32d: color = 2'b10;
      11'h32e: color = 2'b10;
      11'h32f: color = 2'b10;
      11'h330: color = 2'b10;
      11'h331: color = 2'b10;
      11'h332: color = 2'b10;
      11'h333: color = 2'b10;
      11'h334: color = 2'b10;
      11'h335: color = 2'b10;
      11'h336: color = 2'b10;
      11'h337: color = 2'b10;
      11'h338: color = 2'b10;
      11'h339: color = 2'b10;
      11'h33a: color = 2'b00;
      11'h33b: color = 2'b00;
      11'h33c: color = 2'b01;
      11'h33d: color = 2'b01;
      11'h33e: color = 2'b00;
      11'h33f: color = 2'b00;
      11'h340: color = 2'b00;
      11'h341: color = 2'b00;
      11'h342: color = 2'b11;
      11'h343: color = 2'b11;
      11'h344: color = 2'b00;
      11'h345: color = 2'b00;
      11'h346: color = 2'b01;
      11'h347: color = 2'b01;
      11'h348: color = 2'b01;
      11'h349: color = 2'b01;
      11'h34a: color = 2'b01;
      11'h34b: color = 2'b01;
      11'h34c: color = 2'b01;
      11'h34d: color = 2'b01;
      11'h34e: color = 2'b01;
      11'h34f: color = 2'b01;
      11'h350: color = 2'b01;
      11'h351: color = 2'b01;
      11'h352: color = 2'b01;
      11'h353: color = 2'b01;
      11'h354: color = 2'b01;
      11'h355: color = 2'b01;
      11'h356: color = 2'b01;
      11'h357: color = 2'b01;
      11'h358: color = 2'b01;
      11'h359: color = 2'b01;
      11'h35a: color = 2'b00;
      11'h35b: color = 2'b00;
      11'h35c: color = 2'b10;
      11'h35d: color = 2'b10;
      11'h35e: color = 2'b00;
      11'h35f: color = 2'b00;
      11'h360: color = 2'b00;
      11'h361: color = 2'b00;
      11'h362: color = 2'b11;
      11'h363: color = 2'b11;
      11'h364: color = 2'b00;
      11'h365: color = 2'b00;
      11'h366: color = 2'b01;
      11'h367: color = 2'b01;
      11'h368: color = 2'b01;
      11'h369: color = 2'b01;
      11'h36a: color = 2'b01;
      11'h36b: color = 2'b01;
      11'h36c: color = 2'b01;
      11'h36d: color = 2'b01;
      11'h36e: color = 2'b01;
      11'h36f: color = 2'b01;
      11'h370: color = 2'b01;
      11'h371: color = 2'b01;
      11'h372: color = 2'b01;
      11'h373: color = 2'b01;
      11'h374: color = 2'b01;
      11'h375: color = 2'b01;
      11'h376: color = 2'b01;
      11'h377: color = 2'b01;
      11'h378: color = 2'b01;
      11'h379: color = 2'b01;
      11'h37a: color = 2'b00;
      11'h37b: color = 2'b00;
      11'h37c: color = 2'b10;
      11'h37d: color = 2'b10;
      11'h37e: color = 2'b00;
      11'h37f: color = 2'b00;
      11'h380: color = 2'b00;
      11'h381: color = 2'b00;
      11'h382: color = 2'b11;
      11'h383: color = 2'b11;
      11'h384: color = 2'b11;
      11'h385: color = 2'b11;
      11'h386: color = 2'b00;
      11'h387: color = 2'b00;
      11'h388: color = 2'b00;
      11'h389: color = 2'b00;
      11'h38a: color = 2'b00;
      11'h38b: color = 2'b00;
      11'h38c: color = 2'b00;
      11'h38d: color = 2'b00;
      11'h38e: color = 2'b00;
      11'h38f: color = 2'b00;
      11'h390: color = 2'b00;
      11'h391: color = 2'b00;
      11'h392: color = 2'b00;
      11'h393: color = 2'b00;
      11'h394: color = 2'b00;
      11'h395: color = 2'b00;
      11'h396: color = 2'b00;
      11'h397: color = 2'b00;
      11'h398: color = 2'b00;
      11'h399: color = 2'b00;
      11'h39a: color = 2'b10;
      11'h39b: color = 2'b10;
      11'h39c: color = 2'b10;
      11'h39d: color = 2'b10;
      11'h39e: color = 2'b00;
      11'h39f: color = 2'b00;
      11'h3a0: color = 2'b00;
      11'h3a1: color = 2'b00;
      11'h3a2: color = 2'b11;
      11'h3a3: color = 2'b11;
      11'h3a4: color = 2'b11;
      11'h3a5: color = 2'b11;
      11'h3a6: color = 2'b00;
      11'h3a7: color = 2'b00;
      11'h3a8: color = 2'b00;
      11'h3a9: color = 2'b00;
      11'h3aa: color = 2'b00;
      11'h3ab: color = 2'b00;
      11'h3ac: color = 2'b00;
      11'h3ad: color = 2'b00;
      11'h3ae: color = 2'b00;
      11'h3af: color = 2'b00;
      11'h3b0: color = 2'b00;
      11'h3b1: color = 2'b00;
      11'h3b2: color = 2'b00;
      11'h3b3: color = 2'b00;
      11'h3b4: color = 2'b00;
      11'h3b5: color = 2'b00;
      11'h3b6: color = 2'b00;
      11'h3b7: color = 2'b00;
      11'h3b8: color = 2'b00;
      11'h3b9: color = 2'b00;
      11'h3ba: color = 2'b10;
      11'h3bb: color = 2'b10;
      11'h3bc: color = 2'b10;
      11'h3bd: color = 2'b10;
      11'h3be: color = 2'b00;
      11'h3bf: color = 2'b00;
      11'h3c0: color = 2'b00;
      11'h3c1: color = 2'b00;
      11'h3c2: color = 2'b11;
      11'h3c3: color = 2'b11;
      11'h3c4: color = 2'b11;
      11'h3c5: color = 2'b11;
      11'h3c6: color = 2'b11;
      11'h3c7: color = 2'b11;
      11'h3c8: color = 2'b11;
      11'h3c9: color = 2'b11;
      11'h3ca: color = 2'b11;
      11'h3cb: color = 2'b11;
      11'h3cc: color = 2'b11;
      11'h3cd: color = 2'b11;
      11'h3ce: color = 2'b11;
      11'h3cf: color = 2'b11;
      11'h3d0: color = 2'b11;
      11'h3d1: color = 2'b11;
      11'h3d2: color = 2'b11;
      11'h3d3: color = 2'b11;
      11'h3d4: color = 2'b11;
      11'h3d5: color = 2'b11;
      11'h3d6: color = 2'b11;
      11'h3d7: color = 2'b11;
      11'h3d8: color = 2'b11;
      11'h3d9: color = 2'b11;
      11'h3da: color = 2'b11;
      11'h3db: color = 2'b11;
      11'h3dc: color = 2'b11;
      11'h3dd: color = 2'b11;
      11'h3de: color = 2'b00;
      11'h3df: color = 2'b00;
      11'h3e0: color = 2'b00;
      11'h3e1: color = 2'b00;
      11'h3e2: color = 2'b11;
      11'h3e3: color = 2'b11;
      11'h3e4: color = 2'b11;
      11'h3e5: color = 2'b11;
      11'h3e6: color = 2'b11;
      11'h3e7: color = 2'b11;
      11'h3e8: color = 2'b11;
      11'h3e9: color = 2'b11;
      11'h3ea: color = 2'b11;
      11'h3eb: color = 2'b11;
      11'h3ec: color = 2'b11;
      11'h3ed: color = 2'b11;
      11'h3ee: color = 2'b11;
      11'h3ef: color = 2'b11;
      11'h3f0: color = 2'b11;
      11'h3f1: color = 2'b11;
      11'h3f2: color = 2'b11;
      11'h3f3: color = 2'b11;
      11'h3f4: color = 2'b11;
      11'h3f5: color = 2'b11;
      11'h3f6: color = 2'b11;
      11'h3f7: color = 2'b11;
      11'h3f8: color = 2'b11;
      11'h3f9: color = 2'b11;
      11'h3fa: color = 2'b11;
      11'h3fb: color = 2'b11;
      11'h3fc: color = 2'b11;
      11'h3fd: color = 2'b11;
      11'h3fe: color = 2'b00;
      11'h3ff: color = 2'b00;
      11'h400: color = 2'b00;
      11'h401: color = 2'b00;
      11'h402: color = 2'b01;
      11'h403: color = 2'b01;
      11'h404: color = 2'b01;
      11'h405: color = 2'b01;
      11'h406: color = 2'b00;
      11'h407: color = 2'b00;
      11'h408: color = 2'b00;
      11'h409: color = 2'b00;
      11'h40a: color = 2'b00;
      11'h40b: color = 2'b00;
      11'h40c: color = 2'b00;
      11'h40d: color = 2'b00;
      11'h40e: color = 2'b00;
      11'h40f: color = 2'b00;
      11'h410: color = 2'b00;
      11'h411: color = 2'b00;
      11'h412: color = 2'b00;
      11'h413: color = 2'b00;
      11'h414: color = 2'b00;
      11'h415: color = 2'b00;
      11'h416: color = 2'b00;
      11'h417: color = 2'b00;
      11'h418: color = 2'b00;
      11'h419: color = 2'b00;
      11'h41a: color = 2'b01;
      11'h41b: color = 2'b01;
      11'h41c: color = 2'b01;
      11'h41d: color = 2'b01;
      11'h41e: color = 2'b00;
      11'h41f: color = 2'b00;
      11'h420: color = 2'b00;
      11'h421: color = 2'b00;
      11'h422: color = 2'b01;
      11'h423: color = 2'b01;
      11'h424: color = 2'b01;
      11'h425: color = 2'b01;
      11'h426: color = 2'b00;
      11'h427: color = 2'b00;
      11'h428: color = 2'b00;
      11'h429: color = 2'b00;
      11'h42a: color = 2'b00;
      11'h42b: color = 2'b00;
      11'h42c: color = 2'b00;
      11'h42d: color = 2'b00;
      11'h42e: color = 2'b00;
      11'h42f: color = 2'b00;
      11'h430: color = 2'b00;
      11'h431: color = 2'b00;
      11'h432: color = 2'b00;
      11'h433: color = 2'b00;
      11'h434: color = 2'b00;
      11'h435: color = 2'b00;
      11'h436: color = 2'b00;
      11'h437: color = 2'b00;
      11'h438: color = 2'b00;
      11'h439: color = 2'b00;
      11'h43a: color = 2'b01;
      11'h43b: color = 2'b01;
      11'h43c: color = 2'b01;
      11'h43d: color = 2'b01;
      11'h43e: color = 2'b00;
      11'h43f: color = 2'b00;
      11'h440: color = 2'b00;
      11'h441: color = 2'b00;
      11'h442: color = 2'b00;
      11'h443: color = 2'b00;
      11'h444: color = 2'b00;
      11'h445: color = 2'b00;
      11'h446: color = 2'b11;
      11'h447: color = 2'b11;
      11'h448: color = 2'b01;
      11'h449: color = 2'b01;
      11'h44a: color = 2'b11;
      11'h44b: color = 2'b11;
      11'h44c: color = 2'b01;
      11'h44d: color = 2'b01;
      11'h44e: color = 2'b11;
      11'h44f: color = 2'b11;
      11'h450: color = 2'b01;
      11'h451: color = 2'b01;
      11'h452: color = 2'b11;
      11'h453: color = 2'b11;
      11'h454: color = 2'b01;
      11'h455: color = 2'b01;
      11'h456: color = 2'b11;
      11'h457: color = 2'b11;
      11'h458: color = 2'b11;
      11'h459: color = 2'b11;
      11'h45a: color = 2'b00;
      11'h45b: color = 2'b00;
      11'h45c: color = 2'b00;
      11'h45d: color = 2'b00;
      11'h45e: color = 2'b00;
      11'h45f: color = 2'b00;
      11'h460: color = 2'b00;
      11'h461: color = 2'b00;
      11'h462: color = 2'b00;
      11'h463: color = 2'b00;
      11'h464: color = 2'b00;
      11'h465: color = 2'b00;
      11'h466: color = 2'b11;
      11'h467: color = 2'b11;
      11'h468: color = 2'b01;
      11'h469: color = 2'b01;
      11'h46a: color = 2'b11;
      11'h46b: color = 2'b11;
      11'h46c: color = 2'b01;
      11'h46d: color = 2'b01;
      11'h46e: color = 2'b11;
      11'h46f: color = 2'b11;
      11'h470: color = 2'b01;
      11'h471: color = 2'b01;
      11'h472: color = 2'b11;
      11'h473: color = 2'b11;
      11'h474: color = 2'b01;
      11'h475: color = 2'b01;
      11'h476: color = 2'b11;
      11'h477: color = 2'b11;
      11'h478: color = 2'b11;
      11'h479: color = 2'b11;
      11'h47a: color = 2'b00;
      11'h47b: color = 2'b00;
      11'h47c: color = 2'b00;
      11'h47d: color = 2'b00;
      11'h47e: color = 2'b00;
      11'h47f: color = 2'b00;
      11'h480: color = 2'b00;
      11'h481: color = 2'b00;
      11'h482: color = 2'b11;
      11'h483: color = 2'b11;
      11'h484: color = 2'b00;
      11'h485: color = 2'b00;
      11'h486: color = 2'b10;
      11'h487: color = 2'b10;
      11'h488: color = 2'b01;
      11'h489: color = 2'b01;
      11'h48a: color = 2'b01;
      11'h48b: color = 2'b01;
      11'h48c: color = 2'b01;
      11'h48d: color = 2'b01;
      11'h48e: color = 2'b01;
      11'h48f: color = 2'b01;
      11'h490: color = 2'b01;
      11'h491: color = 2'b01;
      11'h492: color = 2'b01;
      11'h493: color = 2'b01;
      11'h494: color = 2'b01;
      11'h495: color = 2'b01;
      11'h496: color = 2'b01;
      11'h497: color = 2'b01;
      11'h498: color = 2'b11;
      11'h499: color = 2'b11;
      11'h49a: color = 2'b00;
      11'h49b: color = 2'b00;
      11'h49c: color = 2'b01;
      11'h49d: color = 2'b01;
      11'h49e: color = 2'b00;
      11'h49f: color = 2'b00;
      11'h4a0: color = 2'b00;
      11'h4a1: color = 2'b00;
      11'h4a2: color = 2'b11;
      11'h4a3: color = 2'b11;
      11'h4a4: color = 2'b00;
      11'h4a5: color = 2'b00;
      11'h4a6: color = 2'b10;
      11'h4a7: color = 2'b10;
      11'h4a8: color = 2'b01;
      11'h4a9: color = 2'b01;
      11'h4aa: color = 2'b01;
      11'h4ab: color = 2'b01;
      11'h4ac: color = 2'b01;
      11'h4ad: color = 2'b01;
      11'h4ae: color = 2'b01;
      11'h4af: color = 2'b01;
      11'h4b0: color = 2'b01;
      11'h4b1: color = 2'b01;
      11'h4b2: color = 2'b01;
      11'h4b3: color = 2'b01;
      11'h4b4: color = 2'b01;
      11'h4b5: color = 2'b01;
      11'h4b6: color = 2'b01;
      11'h4b7: color = 2'b01;
      11'h4b8: color = 2'b11;
      11'h4b9: color = 2'b11;
      11'h4ba: color = 2'b00;
      11'h4bb: color = 2'b00;
      11'h4bc: color = 2'b01;
      11'h4bd: color = 2'b01;
      11'h4be: color = 2'b00;
      11'h4bf: color = 2'b00;
      11'h4c0: color = 2'b00;
      11'h4c1: color = 2'b00;
      11'h4c2: color = 2'b11;
      11'h4c3: color = 2'b11;
      11'h4c4: color = 2'b00;
      11'h4c5: color = 2'b00;
      11'h4c6: color = 2'b11;
      11'h4c7: color = 2'b11;
      11'h4c8: color = 2'b01;
      11'h4c9: color = 2'b01;
      11'h4ca: color = 2'b11;
      11'h4cb: color = 2'b11;
      11'h4cc: color = 2'b01;
      11'h4cd: color = 2'b01;
      11'h4ce: color = 2'b11;
      11'h4cf: color = 2'b11;
      11'h4d0: color = 2'b11;
      11'h4d1: color = 2'b11;
      11'h4d2: color = 2'b11;
      11'h4d3: color = 2'b11;
      11'h4d4: color = 2'b11;
      11'h4d5: color = 2'b11;
      11'h4d6: color = 2'b01;
      11'h4d7: color = 2'b01;
      11'h4d8: color = 2'b11;
      11'h4d9: color = 2'b11;
      11'h4da: color = 2'b00;
      11'h4db: color = 2'b00;
      11'h4dc: color = 2'b01;
      11'h4dd: color = 2'b01;
      11'h4de: color = 2'b00;
      11'h4df: color = 2'b00;
      11'h4e0: color = 2'b00;
      11'h4e1: color = 2'b00;
      11'h4e2: color = 2'b11;
      11'h4e3: color = 2'b11;
      11'h4e4: color = 2'b00;
      11'h4e5: color = 2'b00;
      11'h4e6: color = 2'b11;
      11'h4e7: color = 2'b11;
      11'h4e8: color = 2'b01;
      11'h4e9: color = 2'b01;
      11'h4ea: color = 2'b11;
      11'h4eb: color = 2'b11;
      11'h4ec: color = 2'b01;
      11'h4ed: color = 2'b01;
      11'h4ee: color = 2'b11;
      11'h4ef: color = 2'b11;
      11'h4f0: color = 2'b11;
      11'h4f1: color = 2'b11;
      11'h4f2: color = 2'b11;
      11'h4f3: color = 2'b11;
      11'h4f4: color = 2'b11;
      11'h4f5: color = 2'b11;
      11'h4f6: color = 2'b01;
      11'h4f7: color = 2'b01;
      11'h4f8: color = 2'b11;
      11'h4f9: color = 2'b11;
      11'h4fa: color = 2'b00;
      11'h4fb: color = 2'b00;
      11'h4fc: color = 2'b01;
      11'h4fd: color = 2'b01;
      11'h4fe: color = 2'b00;
      11'h4ff: color = 2'b00;
      11'h500: color = 2'b00;
      11'h501: color = 2'b00;
      11'h502: color = 2'b11;
      11'h503: color = 2'b11;
      11'h504: color = 2'b00;
      11'h505: color = 2'b00;
      11'h506: color = 2'b10;
      11'h507: color = 2'b10;
      11'h508: color = 2'b10;
      11'h509: color = 2'b10;
      11'h50a: color = 2'b10;
      11'h50b: color = 2'b10;
      11'h50c: color = 2'b10;
      11'h50d: color = 2'b10;
      11'h50e: color = 2'b10;
      11'h50f: color = 2'b10;
      11'h510: color = 2'b10;
      11'h511: color = 2'b10;
      11'h512: color = 2'b10;
      11'h513: color = 2'b10;
      11'h514: color = 2'b10;
      11'h515: color = 2'b10;
      11'h516: color = 2'b10;
      11'h517: color = 2'b10;
      11'h518: color = 2'b10;
      11'h519: color = 2'b10;
      11'h51a: color = 2'b00;
      11'h51b: color = 2'b00;
      11'h51c: color = 2'b01;
      11'h51d: color = 2'b01;
      11'h51e: color = 2'b00;
      11'h51f: color = 2'b00;
      11'h520: color = 2'b00;
      11'h521: color = 2'b00;
      11'h522: color = 2'b11;
      11'h523: color = 2'b11;
      11'h524: color = 2'b00;
      11'h525: color = 2'b00;
      11'h526: color = 2'b10;
      11'h527: color = 2'b10;
      11'h528: color = 2'b10;
      11'h529: color = 2'b10;
      11'h52a: color = 2'b10;
      11'h52b: color = 2'b10;
      11'h52c: color = 2'b10;
      11'h52d: color = 2'b10;
      11'h52e: color = 2'b10;
      11'h52f: color = 2'b10;
      11'h530: color = 2'b10;
      11'h531: color = 2'b10;
      11'h532: color = 2'b10;
      11'h533: color = 2'b10;
      11'h534: color = 2'b10;
      11'h535: color = 2'b10;
      11'h536: color = 2'b10;
      11'h537: color = 2'b10;
      11'h538: color = 2'b10;
      11'h539: color = 2'b10;
      11'h53a: color = 2'b00;
      11'h53b: color = 2'b00;
      11'h53c: color = 2'b01;
      11'h53d: color = 2'b01;
      11'h53e: color = 2'b00;
      11'h53f: color = 2'b00;
      11'h540: color = 2'b00;
      11'h541: color = 2'b00;
      11'h542: color = 2'b01;
      11'h543: color = 2'b01;
      11'h544: color = 2'b00;
      11'h545: color = 2'b00;
      11'h546: color = 2'b00;
      11'h547: color = 2'b00;
      11'h548: color = 2'b00;
      11'h549: color = 2'b00;
      11'h54a: color = 2'b00;
      11'h54b: color = 2'b00;
      11'h54c: color = 2'b00;
      11'h54d: color = 2'b00;
      11'h54e: color = 2'b00;
      11'h54f: color = 2'b00;
      11'h550: color = 2'b00;
      11'h551: color = 2'b00;
      11'h552: color = 2'b00;
      11'h553: color = 2'b00;
      11'h554: color = 2'b00;
      11'h555: color = 2'b00;
      11'h556: color = 2'b00;
      11'h557: color = 2'b00;
      11'h558: color = 2'b00;
      11'h559: color = 2'b00;
      11'h55a: color = 2'b00;
      11'h55b: color = 2'b00;
      11'h55c: color = 2'b01;
      11'h55d: color = 2'b01;
      11'h55e: color = 2'b00;
      11'h55f: color = 2'b00;
      11'h560: color = 2'b00;
      11'h561: color = 2'b00;
      11'h562: color = 2'b01;
      11'h563: color = 2'b01;
      11'h564: color = 2'b00;
      11'h565: color = 2'b00;
      11'h566: color = 2'b00;
      11'h567: color = 2'b00;
      11'h568: color = 2'b00;
      11'h569: color = 2'b00;
      11'h56a: color = 2'b00;
      11'h56b: color = 2'b00;
      11'h56c: color = 2'b00;
      11'h56d: color = 2'b00;
      11'h56e: color = 2'b00;
      11'h56f: color = 2'b00;
      11'h570: color = 2'b00;
      11'h571: color = 2'b00;
      11'h572: color = 2'b00;
      11'h573: color = 2'b00;
      11'h574: color = 2'b00;
      11'h575: color = 2'b00;
      11'h576: color = 2'b00;
      11'h577: color = 2'b00;
      11'h578: color = 2'b00;
      11'h579: color = 2'b00;
      11'h57a: color = 2'b00;
      11'h57b: color = 2'b00;
      11'h57c: color = 2'b01;
      11'h57d: color = 2'b01;
      11'h57e: color = 2'b00;
      11'h57f: color = 2'b00;
      11'h580: color = 2'b00;
      11'h581: color = 2'b00;
      11'h582: color = 2'b01;
      11'h583: color = 2'b01;
      11'h584: color = 2'b01;
      11'h585: color = 2'b01;
      11'h586: color = 2'b01;
      11'h587: color = 2'b01;
      11'h588: color = 2'b01;
      11'h589: color = 2'b01;
      11'h58a: color = 2'b01;
      11'h58b: color = 2'b01;
      11'h58c: color = 2'b01;
      11'h58d: color = 2'b01;
      11'h58e: color = 2'b01;
      11'h58f: color = 2'b01;
      11'h590: color = 2'b01;
      11'h591: color = 2'b01;
      11'h592: color = 2'b01;
      11'h593: color = 2'b01;
      11'h594: color = 2'b01;
      11'h595: color = 2'b01;
      11'h596: color = 2'b01;
      11'h597: color = 2'b01;
      11'h598: color = 2'b01;
      11'h599: color = 2'b01;
      11'h59a: color = 2'b01;
      11'h59b: color = 2'b01;
      11'h59c: color = 2'b01;
      11'h59d: color = 2'b01;
      11'h59e: color = 2'b00;
      11'h59f: color = 2'b00;
      11'h5a0: color = 2'b00;
      11'h5a1: color = 2'b00;
      11'h5a2: color = 2'b01;
      11'h5a3: color = 2'b01;
      11'h5a4: color = 2'b01;
      11'h5a5: color = 2'b01;
      11'h5a6: color = 2'b01;
      11'h5a7: color = 2'b01;
      11'h5a8: color = 2'b01;
      11'h5a9: color = 2'b01;
      11'h5aa: color = 2'b01;
      11'h5ab: color = 2'b01;
      11'h5ac: color = 2'b01;
      11'h5ad: color = 2'b01;
      11'h5ae: color = 2'b01;
      11'h5af: color = 2'b01;
      11'h5b0: color = 2'b01;
      11'h5b1: color = 2'b01;
      11'h5b2: color = 2'b01;
      11'h5b3: color = 2'b01;
      11'h5b4: color = 2'b01;
      11'h5b5: color = 2'b01;
      11'h5b6: color = 2'b01;
      11'h5b7: color = 2'b01;
      11'h5b8: color = 2'b01;
      11'h5b9: color = 2'b01;
      11'h5ba: color = 2'b01;
      11'h5bb: color = 2'b01;
      11'h5bc: color = 2'b01;
      11'h5bd: color = 2'b01;
      11'h5be: color = 2'b00;
      11'h5bf: color = 2'b00;
      11'h5c0: color = 2'b11;
      11'h5c1: color = 2'b11;
      11'h5c2: color = 2'b00;
      11'h5c3: color = 2'b00;
      11'h5c4: color = 2'b00;
      11'h5c5: color = 2'b00;
      11'h5c6: color = 2'b00;
      11'h5c7: color = 2'b00;
      11'h5c8: color = 2'b00;
      11'h5c9: color = 2'b00;
      11'h5ca: color = 2'b00;
      11'h5cb: color = 2'b00;
      11'h5cc: color = 2'b00;
      11'h5cd: color = 2'b00;
      11'h5ce: color = 2'b00;
      11'h5cf: color = 2'b00;
      11'h5d0: color = 2'b00;
      11'h5d1: color = 2'b00;
      11'h5d2: color = 2'b00;
      11'h5d3: color = 2'b00;
      11'h5d4: color = 2'b00;
      11'h5d5: color = 2'b00;
      11'h5d6: color = 2'b00;
      11'h5d7: color = 2'b00;
      11'h5d8: color = 2'b00;
      11'h5d9: color = 2'b00;
      11'h5da: color = 2'b00;
      11'h5db: color = 2'b00;
      11'h5dc: color = 2'b00;
      11'h5dd: color = 2'b00;
      11'h5de: color = 2'b11;
      11'h5df: color = 2'b11;
      11'h5e0: color = 2'b11;
      11'h5e1: color = 2'b11;
      11'h5e2: color = 2'b00;
      11'h5e3: color = 2'b00;
      11'h5e4: color = 2'b00;
      11'h5e5: color = 2'b00;
      11'h5e6: color = 2'b00;
      11'h5e7: color = 2'b00;
      11'h5e8: color = 2'b00;
      11'h5e9: color = 2'b00;
      11'h5ea: color = 2'b00;
      11'h5eb: color = 2'b00;
      11'h5ec: color = 2'b00;
      11'h5ed: color = 2'b00;
      11'h5ee: color = 2'b00;
      11'h5ef: color = 2'b00;
      11'h5f0: color = 2'b00;
      11'h5f1: color = 2'b00;
      11'h5f2: color = 2'b00;
      11'h5f3: color = 2'b00;
      11'h5f4: color = 2'b00;
      11'h5f5: color = 2'b00;
      11'h5f6: color = 2'b00;
      11'h5f7: color = 2'b00;
      11'h5f8: color = 2'b00;
      11'h5f9: color = 2'b00;
      11'h5fa: color = 2'b00;
      11'h5fb: color = 2'b00;
      11'h5fc: color = 2'b00;
      11'h5fd: color = 2'b00;
      11'h5fe: color = 2'b11;
      11'h5ff: color = 2'b11;
      11'h600: color = 2'b00;
      11'h601: color = 2'b00;
      11'h602: color = 2'b01;
      11'h603: color = 2'b01;
      11'h604: color = 2'b00;
      11'h605: color = 2'b00;
      11'h606: color = 2'b00;
      11'h607: color = 2'b00;
      11'h608: color = 2'b00;
      11'h609: color = 2'b00;
      11'h60a: color = 2'b00;
      11'h60b: color = 2'b00;
      11'h60c: color = 2'b00;
      11'h60d: color = 2'b00;
      11'h60e: color = 2'b00;
      11'h60f: color = 2'b00;
      11'h610: color = 2'b00;
      11'h611: color = 2'b00;
      11'h612: color = 2'b00;
      11'h613: color = 2'b00;
      11'h614: color = 2'b00;
      11'h615: color = 2'b00;
      11'h616: color = 2'b00;
      11'h617: color = 2'b00;
      11'h618: color = 2'b00;
      11'h619: color = 2'b00;
      11'h61a: color = 2'b00;
      11'h61b: color = 2'b00;
      11'h61c: color = 2'b01;
      11'h61d: color = 2'b01;
      11'h61e: color = 2'b00;
      11'h61f: color = 2'b00;
      11'h620: color = 2'b00;
      11'h621: color = 2'b00;
      11'h622: color = 2'b01;
      11'h623: color = 2'b01;
      11'h624: color = 2'b00;
      11'h625: color = 2'b00;
      11'h626: color = 2'b00;
      11'h627: color = 2'b00;
      11'h628: color = 2'b00;
      11'h629: color = 2'b00;
      11'h62a: color = 2'b00;
      11'h62b: color = 2'b00;
      11'h62c: color = 2'b00;
      11'h62d: color = 2'b00;
      11'h62e: color = 2'b00;
      11'h62f: color = 2'b00;
      11'h630: color = 2'b00;
      11'h631: color = 2'b00;
      11'h632: color = 2'b00;
      11'h633: color = 2'b00;
      11'h634: color = 2'b00;
      11'h635: color = 2'b00;
      11'h636: color = 2'b00;
      11'h637: color = 2'b00;
      11'h638: color = 2'b00;
      11'h639: color = 2'b00;
      11'h63a: color = 2'b00;
      11'h63b: color = 2'b00;
      11'h63c: color = 2'b01;
      11'h63d: color = 2'b01;
      11'h63e: color = 2'b00;
      11'h63f: color = 2'b00;
      11'h640: color = 2'b00;
      11'h641: color = 2'b00;
      11'h642: color = 2'b01;
      11'h643: color = 2'b01;
      11'h644: color = 2'b10;
      11'h645: color = 2'b10;
      11'h646: color = 2'b10;
      11'h647: color = 2'b10;
      11'h648: color = 2'b10;
      11'h649: color = 2'b10;
      11'h64a: color = 2'b10;
      11'h64b: color = 2'b10;
      11'h64c: color = 2'b10;
      11'h64d: color = 2'b10;
      11'h64e: color = 2'b00;
      11'h64f: color = 2'b00;
      11'h650: color = 2'b00;
      11'h651: color = 2'b00;
      11'h652: color = 2'b10;
      11'h653: color = 2'b10;
      11'h654: color = 2'b10;
      11'h655: color = 2'b10;
      11'h656: color = 2'b10;
      11'h657: color = 2'b10;
      11'h658: color = 2'b10;
      11'h659: color = 2'b10;
      11'h65a: color = 2'b10;
      11'h65b: color = 2'b10;
      11'h65c: color = 2'b01;
      11'h65d: color = 2'b01;
      11'h65e: color = 2'b00;
      11'h65f: color = 2'b00;
      11'h660: color = 2'b00;
      11'h661: color = 2'b00;
      11'h662: color = 2'b01;
      11'h663: color = 2'b01;
      11'h664: color = 2'b10;
      11'h665: color = 2'b10;
      11'h666: color = 2'b10;
      11'h667: color = 2'b10;
      11'h668: color = 2'b10;
      11'h669: color = 2'b10;
      11'h66a: color = 2'b10;
      11'h66b: color = 2'b10;
      11'h66c: color = 2'b10;
      11'h66d: color = 2'b10;
      11'h66e: color = 2'b00;
      11'h66f: color = 2'b00;
      11'h670: color = 2'b00;
      11'h671: color = 2'b00;
      11'h672: color = 2'b10;
      11'h673: color = 2'b10;
      11'h674: color = 2'b10;
      11'h675: color = 2'b10;
      11'h676: color = 2'b10;
      11'h677: color = 2'b10;
      11'h678: color = 2'b10;
      11'h679: color = 2'b10;
      11'h67a: color = 2'b10;
      11'h67b: color = 2'b10;
      11'h67c: color = 2'b01;
      11'h67d: color = 2'b01;
      11'h67e: color = 2'b00;
      11'h67f: color = 2'b00;
      11'h680: color = 2'b00;
      11'h681: color = 2'b00;
      11'h682: color = 2'b01;
      11'h683: color = 2'b01;
      11'h684: color = 2'b10;
      11'h685: color = 2'b10;
      11'h686: color = 2'b10;
      11'h687: color = 2'b10;
      11'h688: color = 2'b10;
      11'h689: color = 2'b10;
      11'h68a: color = 2'b10;
      11'h68b: color = 2'b10;
      11'h68c: color = 2'b10;
      11'h68d: color = 2'b10;
      11'h68e: color = 2'b00;
      11'h68f: color = 2'b00;
      11'h690: color = 2'b00;
      11'h691: color = 2'b00;
      11'h692: color = 2'b10;
      11'h693: color = 2'b10;
      11'h694: color = 2'b10;
      11'h695: color = 2'b10;
      11'h696: color = 2'b10;
      11'h697: color = 2'b10;
      11'h698: color = 2'b10;
      11'h699: color = 2'b10;
      11'h69a: color = 2'b10;
      11'h69b: color = 2'b10;
      11'h69c: color = 2'b01;
      11'h69d: color = 2'b01;
      11'h69e: color = 2'b00;
      11'h69f: color = 2'b00;
      11'h6a0: color = 2'b00;
      11'h6a1: color = 2'b00;
      11'h6a2: color = 2'b01;
      11'h6a3: color = 2'b01;
      11'h6a4: color = 2'b10;
      11'h6a5: color = 2'b10;
      11'h6a6: color = 2'b10;
      11'h6a7: color = 2'b10;
      11'h6a8: color = 2'b10;
      11'h6a9: color = 2'b10;
      11'h6aa: color = 2'b10;
      11'h6ab: color = 2'b10;
      11'h6ac: color = 2'b10;
      11'h6ad: color = 2'b10;
      11'h6ae: color = 2'b00;
      11'h6af: color = 2'b00;
      11'h6b0: color = 2'b00;
      11'h6b1: color = 2'b00;
      11'h6b2: color = 2'b10;
      11'h6b3: color = 2'b10;
      11'h6b4: color = 2'b10;
      11'h6b5: color = 2'b10;
      11'h6b6: color = 2'b10;
      11'h6b7: color = 2'b10;
      11'h6b8: color = 2'b10;
      11'h6b9: color = 2'b10;
      11'h6ba: color = 2'b10;
      11'h6bb: color = 2'b10;
      11'h6bc: color = 2'b01;
      11'h6bd: color = 2'b01;
      11'h6be: color = 2'b00;
      11'h6bf: color = 2'b00;
      11'h6c0: color = 2'b00;
      11'h6c1: color = 2'b00;
      11'h6c2: color = 2'b01;
      11'h6c3: color = 2'b01;
      11'h6c4: color = 2'b10;
      11'h6c5: color = 2'b10;
      11'h6c6: color = 2'b10;
      11'h6c7: color = 2'b10;
      11'h6c8: color = 2'b10;
      11'h6c9: color = 2'b10;
      11'h6ca: color = 2'b10;
      11'h6cb: color = 2'b10;
      11'h6cc: color = 2'b10;
      11'h6cd: color = 2'b10;
      11'h6ce: color = 2'b00;
      11'h6cf: color = 2'b00;
      11'h6d0: color = 2'b00;
      11'h6d1: color = 2'b00;
      11'h6d2: color = 2'b10;
      11'h6d3: color = 2'b10;
      11'h6d4: color = 2'b10;
      11'h6d5: color = 2'b10;
      11'h6d6: color = 2'b10;
      11'h6d7: color = 2'b10;
      11'h6d8: color = 2'b10;
      11'h6d9: color = 2'b10;
      11'h6da: color = 2'b10;
      11'h6db: color = 2'b10;
      11'h6dc: color = 2'b01;
      11'h6dd: color = 2'b01;
      11'h6de: color = 2'b00;
      11'h6df: color = 2'b00;
      11'h6e0: color = 2'b00;
      11'h6e1: color = 2'b00;
      11'h6e2: color = 2'b01;
      11'h6e3: color = 2'b01;
      11'h6e4: color = 2'b10;
      11'h6e5: color = 2'b10;
      11'h6e6: color = 2'b10;
      11'h6e7: color = 2'b10;
      11'h6e8: color = 2'b10;
      11'h6e9: color = 2'b10;
      11'h6ea: color = 2'b10;
      11'h6eb: color = 2'b10;
      11'h6ec: color = 2'b10;
      11'h6ed: color = 2'b10;
      11'h6ee: color = 2'b00;
      11'h6ef: color = 2'b00;
      11'h6f0: color = 2'b00;
      11'h6f1: color = 2'b00;
      11'h6f2: color = 2'b10;
      11'h6f3: color = 2'b10;
      11'h6f4: color = 2'b10;
      11'h6f5: color = 2'b10;
      11'h6f6: color = 2'b10;
      11'h6f7: color = 2'b10;
      11'h6f8: color = 2'b10;
      11'h6f9: color = 2'b10;
      11'h6fa: color = 2'b10;
      11'h6fb: color = 2'b10;
      11'h6fc: color = 2'b01;
      11'h6fd: color = 2'b01;
      11'h6fe: color = 2'b00;
      11'h6ff: color = 2'b00;
      11'h700: color = 2'b00;
      11'h701: color = 2'b00;
      11'h702: color = 2'b01;
      11'h703: color = 2'b01;
      11'h704: color = 2'b10;
      11'h705: color = 2'b10;
      11'h706: color = 2'b10;
      11'h707: color = 2'b10;
      11'h708: color = 2'b10;
      11'h709: color = 2'b10;
      11'h70a: color = 2'b10;
      11'h70b: color = 2'b10;
      11'h70c: color = 2'b10;
      11'h70d: color = 2'b10;
      11'h70e: color = 2'b00;
      11'h70f: color = 2'b00;
      11'h710: color = 2'b00;
      11'h711: color = 2'b00;
      11'h712: color = 2'b10;
      11'h713: color = 2'b10;
      11'h714: color = 2'b10;
      11'h715: color = 2'b10;
      11'h716: color = 2'b10;
      11'h717: color = 2'b10;
      11'h718: color = 2'b10;
      11'h719: color = 2'b10;
      11'h71a: color = 2'b10;
      11'h71b: color = 2'b10;
      11'h71c: color = 2'b01;
      11'h71d: color = 2'b01;
      11'h71e: color = 2'b00;
      11'h71f: color = 2'b00;
      11'h720: color = 2'b00;
      11'h721: color = 2'b00;
      11'h722: color = 2'b01;
      11'h723: color = 2'b01;
      11'h724: color = 2'b10;
      11'h725: color = 2'b10;
      11'h726: color = 2'b10;
      11'h727: color = 2'b10;
      11'h728: color = 2'b10;
      11'h729: color = 2'b10;
      11'h72a: color = 2'b10;
      11'h72b: color = 2'b10;
      11'h72c: color = 2'b10;
      11'h72d: color = 2'b10;
      11'h72e: color = 2'b00;
      11'h72f: color = 2'b00;
      11'h730: color = 2'b00;
      11'h731: color = 2'b00;
      11'h732: color = 2'b10;
      11'h733: color = 2'b10;
      11'h734: color = 2'b10;
      11'h735: color = 2'b10;
      11'h736: color = 2'b10;
      11'h737: color = 2'b10;
      11'h738: color = 2'b10;
      11'h739: color = 2'b10;
      11'h73a: color = 2'b10;
      11'h73b: color = 2'b10;
      11'h73c: color = 2'b01;
      11'h73d: color = 2'b01;
      11'h73e: color = 2'b00;
      11'h73f: color = 2'b00;
      11'h740: color = 2'b00;
      11'h741: color = 2'b00;
      11'h742: color = 2'b00;
      11'h743: color = 2'b00;
      11'h744: color = 2'b00;
      11'h745: color = 2'b00;
      11'h746: color = 2'b00;
      11'h747: color = 2'b00;
      11'h748: color = 2'b00;
      11'h749: color = 2'b00;
      11'h74a: color = 2'b00;
      11'h74b: color = 2'b00;
      11'h74c: color = 2'b00;
      11'h74d: color = 2'b00;
      11'h74e: color = 2'b00;
      11'h74f: color = 2'b00;
      11'h750: color = 2'b00;
      11'h751: color = 2'b00;
      11'h752: color = 2'b00;
      11'h753: color = 2'b00;
      11'h754: color = 2'b00;
      11'h755: color = 2'b00;
      11'h756: color = 2'b00;
      11'h757: color = 2'b00;
      11'h758: color = 2'b00;
      11'h759: color = 2'b00;
      11'h75a: color = 2'b00;
      11'h75b: color = 2'b00;
      11'h75c: color = 2'b00;
      11'h75d: color = 2'b00;
      11'h75e: color = 2'b00;
      11'h75f: color = 2'b00;
      11'h760: color = 2'b00;
      11'h761: color = 2'b00;
      11'h762: color = 2'b00;
      11'h763: color = 2'b00;
      11'h764: color = 2'b00;
      11'h765: color = 2'b00;
      11'h766: color = 2'b00;
      11'h767: color = 2'b00;
      11'h768: color = 2'b00;
      11'h769: color = 2'b00;
      11'h76a: color = 2'b00;
      11'h76b: color = 2'b00;
      11'h76c: color = 2'b00;
      11'h76d: color = 2'b00;
      11'h76e: color = 2'b00;
      11'h76f: color = 2'b00;
      11'h770: color = 2'b00;
      11'h771: color = 2'b00;
      11'h772: color = 2'b00;
      11'h773: color = 2'b00;
      11'h774: color = 2'b00;
      11'h775: color = 2'b00;
      11'h776: color = 2'b00;
      11'h777: color = 2'b00;
      11'h778: color = 2'b00;
      11'h779: color = 2'b00;
      11'h77a: color = 2'b00;
      11'h77b: color = 2'b00;
      11'h77c: color = 2'b00;
      11'h77d: color = 2'b00;
      11'h77e: color = 2'b00;
      11'h77f: color = 2'b00;
      11'h780: color = 2'b00;
      11'h781: color = 2'b00;
      11'h782: color = 2'b01;
      11'h783: color = 2'b01;
      11'h784: color = 2'b10;
      11'h785: color = 2'b10;
      11'h786: color = 2'b10;
      11'h787: color = 2'b10;
      11'h788: color = 2'b10;
      11'h789: color = 2'b10;
      11'h78a: color = 2'b10;
      11'h78b: color = 2'b10;
      11'h78c: color = 2'b10;
      11'h78d: color = 2'b10;
      11'h78e: color = 2'b10;
      11'h78f: color = 2'b10;
      11'h790: color = 2'b10;
      11'h791: color = 2'b10;
      11'h792: color = 2'b10;
      11'h793: color = 2'b10;
      11'h794: color = 2'b10;
      11'h795: color = 2'b10;
      11'h796: color = 2'b10;
      11'h797: color = 2'b10;
      11'h798: color = 2'b10;
      11'h799: color = 2'b10;
      11'h79a: color = 2'b10;
      11'h79b: color = 2'b10;
      11'h79c: color = 2'b01;
      11'h79d: color = 2'b01;
      11'h79e: color = 2'b00;
      11'h79f: color = 2'b00;
      11'h7a0: color = 2'b00;
      11'h7a1: color = 2'b00;
      11'h7a2: color = 2'b01;
      11'h7a3: color = 2'b01;
      11'h7a4: color = 2'b10;
      11'h7a5: color = 2'b10;
      11'h7a6: color = 2'b10;
      11'h7a7: color = 2'b10;
      11'h7a8: color = 2'b10;
      11'h7a9: color = 2'b10;
      11'h7aa: color = 2'b10;
      11'h7ab: color = 2'b10;
      11'h7ac: color = 2'b10;
      11'h7ad: color = 2'b10;
      11'h7ae: color = 2'b10;
      11'h7af: color = 2'b10;
      11'h7b0: color = 2'b10;
      11'h7b1: color = 2'b10;
      11'h7b2: color = 2'b10;
      11'h7b3: color = 2'b10;
      11'h7b4: color = 2'b10;
      11'h7b5: color = 2'b10;
      11'h7b6: color = 2'b10;
      11'h7b7: color = 2'b10;
      11'h7b8: color = 2'b10;
      11'h7b9: color = 2'b10;
      11'h7ba: color = 2'b10;
      11'h7bb: color = 2'b10;
      11'h7bc: color = 2'b01;
      11'h7bd: color = 2'b01;
      11'h7be: color = 2'b00;
      11'h7bf: color = 2'b00;
      11'h7c0: color = 2'b11;
      11'h7c1: color = 2'b11;
      11'h7c2: color = 2'b00;
      11'h7c3: color = 2'b00;
      11'h7c4: color = 2'b00;
      11'h7c5: color = 2'b00;
      11'h7c6: color = 2'b00;
      11'h7c7: color = 2'b00;
      11'h7c8: color = 2'b00;
      11'h7c9: color = 2'b00;
      11'h7ca: color = 2'b00;
      11'h7cb: color = 2'b00;
      11'h7cc: color = 2'b00;
      11'h7cd: color = 2'b00;
      11'h7ce: color = 2'b00;
      11'h7cf: color = 2'b00;
      11'h7d0: color = 2'b00;
      11'h7d1: color = 2'b00;
      11'h7d2: color = 2'b00;
      11'h7d3: color = 2'b00;
      11'h7d4: color = 2'b00;
      11'h7d5: color = 2'b00;
      11'h7d6: color = 2'b00;
      11'h7d7: color = 2'b00;
      11'h7d8: color = 2'b00;
      11'h7d9: color = 2'b00;
      11'h7da: color = 2'b00;
      11'h7db: color = 2'b00;
      11'h7dc: color = 2'b00;
      11'h7dd: color = 2'b00;
      11'h7de: color = 2'b11;
      11'h7df: color = 2'b11;
      11'h7e0: color = 2'b11;
      11'h7e1: color = 2'b11;
      11'h7e2: color = 2'b00;
      11'h7e3: color = 2'b00;
      11'h7e4: color = 2'b00;
      11'h7e5: color = 2'b00;
      11'h7e6: color = 2'b00;
      11'h7e7: color = 2'b00;
      11'h7e8: color = 2'b00;
      11'h7e9: color = 2'b00;
      11'h7ea: color = 2'b00;
      11'h7eb: color = 2'b00;
      11'h7ec: color = 2'b00;
      11'h7ed: color = 2'b00;
      11'h7ee: color = 2'b00;
      11'h7ef: color = 2'b00;
      11'h7f0: color = 2'b00;
      11'h7f1: color = 2'b00;
      11'h7f2: color = 2'b00;
      11'h7f3: color = 2'b00;
      11'h7f4: color = 2'b00;
      11'h7f5: color = 2'b00;
      11'h7f6: color = 2'b00;
      11'h7f7: color = 2'b00;
      11'h7f8: color = 2'b00;
      11'h7f9: color = 2'b00;
      11'h7fa: color = 2'b00;
      11'h7fb: color = 2'b00;
      11'h7fc: color = 2'b00;
      11'h7fd: color = 2'b00;
      11'h7fe: color = 2'b11;
      11'h7ff: color = 2'b11;
      default: color = 2'b11;
   endcase
end
endmodule
